library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity bpsk_modulator is
    Port ( clk : in STD_LOGIC;
           tx : in STD_LOGIC;
           baseband : out STD_LOGIC_VECTOR (15 downto 0));
end bpsk_modulator;

architecture Behavioral of bpsk_modulator is
   type a_lookup is array(0 to 8191) of std_logic_vector(15 downto 0);
   signal lookup : a_lookup := (
        x"92a1", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0",
        x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0", x"92a0",
        x"92a0", x"92a0", x"92a0", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f",
        x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f", x"929f",
        x"929f", x"929f", x"929f", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e",
        x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e", x"929e",
        x"929e", x"929e", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d",
        x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929d", x"929c",
        x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c",
        x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929c", x"929b", x"929b", x"929b", x"929b", x"929b", x"929b", x"929b",
        x"929b", x"929b", x"929b", x"929b", x"929b", x"929b", x"929b", x"929b", x"929b", x"929b", x"929b", x"929b", x"929b", x"929b", x"929b", x"929b",
        x"929b", x"929b", x"929b", x"929a", x"929a", x"929a", x"929a", x"929a", x"929a", x"929a", x"929a", x"929a", x"929a", x"929a", x"929a", x"929a",
        x"929a", x"929a", x"929a", x"929a", x"929a", x"929a", x"929a", x"929a", x"929a", x"929a", x"9299", x"9299", x"9299", x"9299", x"9299", x"9299",
        x"9299", x"9299", x"9299", x"9299", x"9299", x"9299", x"9299", x"9299", x"9299", x"9299", x"9299", x"9299", x"9299", x"9299", x"9299", x"9299",
        x"9298", x"9298", x"9298", x"9298", x"9298", x"9298", x"9298", x"9298", x"9298", x"9298", x"9298", x"9298", x"9298", x"9298", x"9298", x"9298",
        x"9298", x"9298", x"9298", x"9298", x"9297", x"9297", x"9297", x"9297", x"9297", x"9297", x"9297", x"9297", x"9297", x"9297", x"9297", x"9297",
        x"9297", x"9297", x"9297", x"9297", x"9297", x"9297", x"9297", x"9297", x"9296", x"9296", x"9296", x"9296", x"9296", x"9296", x"9296", x"9296",
        x"9296", x"9296", x"9296", x"9296", x"9296", x"9296", x"9296", x"9296", x"9296", x"9296", x"9295", x"9295", x"9295", x"9295", x"9295", x"9295",
        x"9295", x"9295", x"9295", x"9295", x"9295", x"9295", x"9295", x"9295", x"9295", x"9295", x"9295", x"9294", x"9294", x"9294", x"9294", x"9294",
        x"9294", x"9294", x"9294", x"9294", x"9294", x"9294", x"9294", x"9294", x"9294", x"9294", x"9294", x"9293", x"9293", x"9293", x"9293", x"9293",
        x"9293", x"9293", x"9293", x"9293", x"9293", x"9293", x"9293", x"9293", x"9293", x"9293", x"9293", x"9292", x"9292", x"9292", x"9292", x"9292",
        x"9292", x"9292", x"9292", x"9292", x"9292", x"9292", x"9292", x"9292", x"9292", x"9292", x"9291", x"9291", x"9291", x"9291", x"9291", x"9291",
        x"9291", x"9291", x"9291", x"9291", x"9291", x"9291", x"9291", x"9291", x"9290", x"9290", x"9290", x"9290", x"9290", x"9290", x"9290", x"9290",
        x"9290", x"9290", x"9290", x"9290", x"9290", x"928f", x"928f", x"928f", x"928f", x"928f", x"928f", x"928f", x"928f", x"928f", x"928f", x"928f",
        x"928f", x"928f", x"928e", x"928e", x"928e", x"928e", x"928e", x"928e", x"928e", x"928e", x"928e", x"928e", x"928e", x"928e", x"928d", x"928d",
        x"928d", x"928d", x"928d", x"928d", x"928d", x"928d", x"928d", x"928d", x"928d", x"928d", x"928c", x"928c", x"928c", x"928c", x"928c", x"928c",
        x"928c", x"928c", x"928c", x"928c", x"928c", x"928c", x"928b", x"928b", x"928b", x"928b", x"928b", x"928b", x"928b", x"928b", x"928b", x"928b",
        x"928b", x"928a", x"928a", x"928a", x"928a", x"928a", x"928a", x"928a", x"928a", x"928a", x"928a", x"928a", x"9289", x"9289", x"9289", x"9289",
        x"9289", x"9289", x"9289", x"9289", x"9289", x"9289", x"9288", x"9288", x"9288", x"9288", x"9288", x"9288", x"9288", x"9288", x"9288", x"9288",
        x"9287", x"9287", x"9287", x"9287", x"9287", x"9287", x"9287", x"9287", x"9287", x"9287", x"9286", x"9286", x"9286", x"9286", x"9286", x"9286",
        x"9286", x"9286", x"9286", x"9286", x"9285", x"9285", x"9285", x"9285", x"9285", x"9285", x"9285", x"9285", x"9285", x"9284", x"9284", x"9284",
        x"9284", x"9284", x"9284", x"9284", x"9284", x"9284", x"9283", x"9283", x"9283", x"9283", x"9283", x"9283", x"9283", x"9283", x"9283", x"9282",
        x"9282", x"9282", x"9282", x"9282", x"9282", x"9282", x"9282", x"9281", x"9281", x"9281", x"9281", x"9281", x"9281", x"9281", x"9281", x"9281",
        x"9280", x"9280", x"9280", x"9280", x"9280", x"9280", x"9280", x"9280", x"927f", x"927f", x"927f", x"927f", x"927f", x"927f", x"927f", x"927f",
        x"927e", x"927e", x"927e", x"927e", x"927e", x"927e", x"927e", x"927e", x"927d", x"927d", x"927d", x"927d", x"927d", x"927d", x"927d", x"927c",
        x"927c", x"927c", x"927c", x"927c", x"927c", x"927c", x"927c", x"927b", x"927b", x"927b", x"927b", x"927b", x"927b", x"927b", x"927a", x"927a",
        x"927a", x"927a", x"927a", x"927a", x"927a", x"927a", x"9279", x"9279", x"9279", x"9279", x"9279", x"9279", x"9279", x"9278", x"9278", x"9278",
        x"9278", x"9278", x"9278", x"9278", x"9277", x"9277", x"9277", x"9277", x"9277", x"9277", x"9277", x"9276", x"9276", x"9276", x"9276", x"9276",
        x"9276", x"9275", x"9275", x"9275", x"9275", x"9275", x"9275", x"9275", x"9274", x"9274", x"9274", x"9274", x"9274", x"9274", x"9273", x"9273",
        x"9273", x"9273", x"9273", x"9273", x"9273", x"9272", x"9272", x"9272", x"9272", x"9272", x"9272", x"9271", x"9271", x"9271", x"9271", x"9271",
        x"9271", x"9270", x"9270", x"9270", x"9270", x"9270", x"9270", x"9270", x"926f", x"926f", x"926f", x"926f", x"926f", x"926f", x"926e", x"926e",
        x"926e", x"926e", x"926e", x"926e", x"926d", x"926d", x"926d", x"926d", x"926d", x"926c", x"926c", x"926c", x"926c", x"926c", x"926c", x"926b",
        x"926b", x"926b", x"926b", x"926b", x"926b", x"926a", x"926a", x"926a", x"926a", x"926a", x"926a", x"9269", x"9269", x"9269", x"9269", x"9269",
        x"9268", x"9268", x"9268", x"9268", x"9268", x"9268", x"9267", x"9267", x"9267", x"9267", x"9267", x"9266", x"9266", x"9266", x"9266", x"9266",
        x"9265", x"9265", x"9265", x"9265", x"9265", x"9265", x"9264", x"9264", x"9264", x"9264", x"9264", x"9263", x"9263", x"9263", x"9263", x"9263",
        x"9262", x"9262", x"9262", x"9262", x"9262", x"9261", x"9261", x"9261", x"9261", x"9261", x"9260", x"9260", x"9260", x"9260", x"9260", x"925f",
        x"925f", x"925f", x"925f", x"925f", x"925e", x"925e", x"925e", x"925e", x"925e", x"925d", x"925d", x"925d", x"925d", x"925d", x"925c", x"925c",
        x"925c", x"925c", x"925c", x"925b", x"925b", x"925b", x"925b", x"925b", x"925a", x"925a", x"925a", x"925a", x"925a", x"9259", x"9259", x"9259",
        x"9259", x"9258", x"9258", x"9258", x"9258", x"9258", x"9257", x"9257", x"9257", x"9257", x"9257", x"9256", x"9256", x"9256", x"9256", x"9255",
        x"9255", x"9255", x"9255", x"9255", x"9254", x"9254", x"9254", x"9254", x"9253", x"9253", x"9253", x"9253", x"9253", x"9252", x"9252", x"9252",
        x"9252", x"9251", x"9251", x"9251", x"9251", x"9250", x"9250", x"9250", x"9250", x"9250", x"924f", x"924f", x"924f", x"924f", x"924e", x"924e",
        x"924e", x"924e", x"924d", x"924d", x"924d", x"924d", x"924d", x"924c", x"924c", x"924c", x"924c", x"924b", x"924b", x"924b", x"924b", x"924a",
        x"924a", x"924a", x"924a", x"9249", x"9249", x"9249", x"9249", x"9248", x"9248", x"9248", x"9248", x"9248", x"9247", x"9247", x"9247", x"9247",
        x"9246", x"9246", x"9246", x"9246", x"9245", x"9245", x"9245", x"9245", x"9244", x"9244", x"9244", x"9244", x"9243", x"9243", x"9243", x"9243",
        x"9242", x"9242", x"9242", x"9242", x"9241", x"9241", x"9241", x"9241", x"9240", x"9240", x"9240", x"923f", x"923f", x"923f", x"923f", x"923e",
        x"923e", x"923e", x"923e", x"923d", x"923d", x"923d", x"923d", x"923c", x"923c", x"923c", x"923c", x"923b", x"923b", x"923b", x"923b", x"923a",
        x"923a", x"923a", x"9239", x"9239", x"9239", x"9239", x"9238", x"9238", x"9238", x"9238", x"9237", x"9237", x"9237", x"9237", x"9236", x"9236",
        x"9236", x"9235", x"9235", x"9235", x"9235", x"9234", x"9234", x"9234", x"9234", x"9233", x"9233", x"9233", x"9232", x"9232", x"9232", x"9232",
        x"9231", x"9231", x"9231", x"9230", x"9230", x"9230", x"9230", x"922f", x"922f", x"922f", x"922f", x"922e", x"922e", x"922e", x"922d", x"922d",
        x"922d", x"922d", x"922c", x"922c", x"922c", x"922b", x"922b", x"922b", x"922b", x"922a", x"922a", x"922a", x"9229", x"9229", x"9229", x"9229",
        x"9228", x"9228", x"9228", x"9227", x"9227", x"9227", x"9226", x"9226", x"9226", x"9226", x"9225", x"9225", x"9225", x"9224", x"9224", x"9224",
        x"9224", x"9223", x"9223", x"9223", x"9222", x"9222", x"9222", x"9221", x"9221", x"9221", x"9221", x"9220", x"9220", x"9220", x"921f", x"921f",
        x"921f", x"921f", x"921e", x"921e", x"921e", x"921d", x"921d", x"921d", x"921c", x"921c", x"921c", x"921c", x"921b", x"921b", x"921b", x"921a",
        x"921a", x"921a", x"9219", x"9219", x"9219", x"9218", x"9218", x"9218", x"9218", x"9217", x"9217", x"9217", x"9216", x"9216", x"9216", x"9215",
        x"9215", x"9215", x"9214", x"9214", x"9214", x"9214", x"9213", x"9213", x"9213", x"9212", x"9212", x"9212", x"9211", x"9211", x"9211", x"9210",
        x"9210", x"9210", x"920f", x"920f", x"920f", x"920f", x"920e", x"920e", x"920e", x"920d", x"920d", x"920d", x"920c", x"920c", x"920c", x"920b",
        x"920b", x"920b", x"920a", x"920a", x"920a", x"9209", x"9209", x"9209", x"9209", x"9208", x"9208", x"9208", x"9207", x"9207", x"9207", x"9206",
        x"9206", x"9206", x"9205", x"9205", x"9205", x"9204", x"9204", x"9204", x"9203", x"9203", x"9203", x"9202", x"9202", x"9202", x"9201", x"9201",
        x"9201", x"9200", x"9200", x"9200", x"9200", x"91ff", x"91ff", x"91ff", x"91fe", x"91fe", x"91fe", x"91fd", x"91fd", x"91fd", x"91fc", x"91fc",
        x"91fc", x"91fb", x"91fb", x"91fb", x"91fa", x"91fa", x"91fa", x"91f9", x"91f9", x"91f9", x"91f8", x"91f8", x"91f8", x"91f7", x"91f7", x"91f7",
        x"91f6", x"91f6", x"91f6", x"91f5", x"91f5", x"91f5", x"91f4", x"91f4", x"91f4", x"91f3", x"91f3", x"91f3", x"91f2", x"91f2", x"91f2", x"91f1",
        x"91f1", x"91f1", x"91f0", x"91f0", x"91f0", x"91ef", x"91ef", x"91ef", x"91ee", x"91ee", x"91ee", x"91ed", x"91ed", x"91ed", x"91ec", x"91ec",
        x"91ec", x"91eb", x"91eb", x"91eb", x"91ea", x"91ea", x"91ea", x"91e9", x"91e9", x"91e9", x"91e8", x"91e8", x"91e8", x"91e7", x"91e7", x"91e7",
        x"91e6", x"91e6", x"91e6", x"91e5", x"91e5", x"91e5", x"91e4", x"91e4", x"91e4", x"91e3", x"91e3", x"91e3", x"91e2", x"91e2", x"91e2", x"91e1",
        x"91e1", x"91e1", x"91e0", x"91e0", x"91e0", x"91df", x"91df", x"91df", x"91de", x"91de", x"91de", x"91dd", x"91dd", x"91dd", x"91dd", x"91dc",
        x"91dc", x"91dc", x"91db", x"91db", x"91db", x"91da", x"91da", x"91da", x"91d9", x"91d9", x"91d9", x"91d8", x"91d8", x"91d8", x"91d7", x"91d7",
        x"91d7", x"91d6", x"91d6", x"91d6", x"91d5", x"91d5", x"91d5", x"91d4", x"91d4", x"91d4", x"91d3", x"91d3", x"91d3", x"91d2", x"91d2", x"91d2",
        x"91d1", x"91d1", x"91d1", x"91d0", x"91d0", x"91d0", x"91cf", x"91cf", x"91cf", x"91ce", x"91ce", x"91ce", x"91cd", x"91cd", x"91cd", x"91cc",
        x"91cc", x"91cc", x"91cb", x"91cb", x"91cb", x"91ca", x"91ca", x"91ca", x"91c9", x"91c9", x"91c9", x"91c8", x"91c8", x"91c8", x"91c7", x"91c7",
        x"91c7", x"91c7", x"91c6", x"91c6", x"91c6", x"91c5", x"91c5", x"91c5", x"91c4", x"91c4", x"91c4", x"91c3", x"91c3", x"91c3", x"91c2", x"91c2",
        x"91c2", x"91c1", x"91c1", x"91c1", x"91c0", x"91c0", x"91c0", x"91bf", x"91bf", x"91bf", x"91bf", x"91be", x"91be", x"91be", x"91bd", x"91bd",
        x"91bd", x"91bc", x"91bc", x"91bc", x"91bb", x"91bb", x"91bb", x"91ba", x"91ba", x"91ba", x"91ba", x"91b9", x"91b9", x"91b9", x"91b8", x"91b8",
        x"91b8", x"91b7", x"91b7", x"91b7", x"91b6", x"91b6", x"91b6", x"91b6", x"91b5", x"91b5", x"91b5", x"91b4", x"91b4", x"91b4", x"91b3", x"91b3",
        x"91b3", x"91b3", x"91b2", x"91b2", x"91b2", x"91b1", x"91b1", x"91b1", x"91b0", x"91b0", x"91b0", x"91b0", x"91af", x"91af", x"91af", x"91ae",
        x"91ae", x"91ae", x"91ae", x"91ad", x"91ad", x"91ad", x"91ac", x"91ac", x"91ac", x"91ac", x"91ab", x"91ab", x"91ab", x"91aa", x"91aa", x"91aa",
        x"91aa", x"91a9", x"91a9", x"91a9", x"91a8", x"91a8", x"91a8", x"91a8", x"91a7", x"91a7", x"91a7", x"91a6", x"91a6", x"91a6", x"91a6", x"91a5",
        x"91a5", x"91a5", x"91a5", x"91a4", x"91a4", x"91a4", x"91a3", x"91a3", x"91a3", x"91a3", x"91a2", x"91a2", x"91a2", x"91a2", x"91a1", x"91a1",
        x"91a1", x"91a1", x"91a0", x"91a0", x"91a0", x"919f", x"919f", x"919f", x"919f", x"919e", x"919e", x"919e", x"919e", x"919d", x"919d", x"919d",
        x"919d", x"919c", x"919c", x"919c", x"919c", x"919b", x"919b", x"919b", x"919b", x"919a", x"919a", x"919a", x"919a", x"919a", x"9199", x"9199",
        x"9199", x"9199", x"9198", x"9198", x"9198", x"9198", x"9197", x"9197", x"9197", x"9197", x"9197", x"9196", x"9196", x"9196", x"9196", x"9195",
        x"9195", x"9195", x"9195", x"9195", x"9194", x"9194", x"9194", x"9194", x"9193", x"9193", x"9193", x"9193", x"9193", x"9192", x"9192", x"9192",
        x"9192", x"9192", x"9191", x"9191", x"9191", x"9191", x"9191", x"9190", x"9190", x"9190", x"9190", x"9190", x"918f", x"918f", x"918f", x"918f",
        x"918f", x"918e", x"918e", x"918e", x"918e", x"918e", x"918e", x"918d", x"918d", x"918d", x"918d", x"918d", x"918c", x"918c", x"918c", x"918c",
        x"918c", x"918c", x"918b", x"918b", x"918b", x"918b", x"918b", x"918b", x"918a", x"918a", x"918a", x"918a", x"918a", x"918a", x"918a", x"9189",
        x"9189", x"9189", x"9189", x"9189", x"9189", x"9189", x"9188", x"9188", x"9188", x"9188", x"9188", x"9188", x"9188", x"9187", x"9187", x"9187",
        x"9187", x"9187", x"9187", x"9187", x"9187", x"9186", x"9186", x"9186", x"9186", x"9186", x"9186", x"9186", x"9186", x"9186", x"9185", x"9185",
        x"9185", x"9185", x"9185", x"9185", x"9185", x"9185", x"9185", x"9185", x"9184", x"9184", x"9184", x"9184", x"9184", x"9184", x"9184", x"9184",
        x"9184", x"9184", x"9184", x"9184", x"9184", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183",
        x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182",
        x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182",
        x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182", x"9182",
        x"9182", x"9182", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183", x"9183",
        x"9183", x"9183", x"9183", x"9184", x"9184", x"9184", x"9184", x"9184", x"9184", x"9184", x"9184", x"9184", x"9184", x"9184", x"9185", x"9185",
        x"9185", x"9185", x"9185", x"9185", x"9185", x"9185", x"9185", x"9186", x"9186", x"9186", x"9186", x"9186", x"9186", x"9186", x"9187", x"9187",
        x"9187", x"9187", x"9187", x"9187", x"9187", x"9188", x"9188", x"9188", x"9188", x"9188", x"9188", x"9189", x"9189", x"9189", x"9189", x"9189",
        x"9189", x"918a", x"918a", x"918a", x"918a", x"918a", x"918b", x"918b", x"918b", x"918b", x"918b", x"918c", x"918c", x"918c", x"918c", x"918d",
        x"918d", x"918d", x"918d", x"918e", x"918e", x"918e", x"918e", x"918e", x"918f", x"918f", x"918f", x"918f", x"9190", x"9190", x"9190", x"9191",
        x"9191", x"9191", x"9191", x"9192", x"9192", x"9192", x"9192", x"9193", x"9193", x"9193", x"9194", x"9194", x"9194", x"9195", x"9195", x"9195",
        x"9195", x"9196", x"9196", x"9196", x"9197", x"9197", x"9197", x"9198", x"9198", x"9198", x"9199", x"9199", x"919a", x"919a", x"919a", x"919b",
        x"919b", x"919b", x"919c", x"919c", x"919c", x"919d", x"919d", x"919e", x"919e", x"919e", x"919f", x"919f", x"91a0", x"91a0", x"91a0", x"91a1",
        x"91a1", x"91a2", x"91a2", x"91a2", x"91a3", x"91a3", x"91a4", x"91a4", x"91a5", x"91a5", x"91a6", x"91a6", x"91a6", x"91a7", x"91a7", x"91a8",
        x"91a8", x"91a9", x"91a9", x"91aa", x"91aa", x"91ab", x"91ab", x"91ac", x"91ac", x"91ad", x"91ad", x"91ae", x"91ae", x"91af", x"91af", x"91b0",
        x"91b0", x"91b1", x"91b1", x"91b2", x"91b2", x"91b3", x"91b3", x"91b4", x"91b4", x"91b5", x"91b6", x"91b6", x"91b7", x"91b7", x"91b8", x"91b8",
        x"91b9", x"91ba", x"91ba", x"91bb", x"91bb", x"91bc", x"91bd", x"91bd", x"91be", x"91be", x"91bf", x"91c0", x"91c0", x"91c1", x"91c1", x"91c2",
        x"91c3", x"91c3", x"91c4", x"91c5", x"91c5", x"91c6", x"91c7", x"91c7", x"91c8", x"91c9", x"91c9", x"91ca", x"91cb", x"91cb", x"91cc", x"91cd",
        x"91cd", x"91ce", x"91cf", x"91d0", x"91d0", x"91d1", x"91d2", x"91d3", x"91d3", x"91d4", x"91d5", x"91d5", x"91d6", x"91d7", x"91d8", x"91d8",
        x"91d9", x"91da", x"91db", x"91dc", x"91dc", x"91dd", x"91de", x"91df", x"91e0", x"91e0", x"91e1", x"91e2", x"91e3", x"91e4", x"91e4", x"91e5",
        x"91e6", x"91e7", x"91e8", x"91e9", x"91e9", x"91ea", x"91eb", x"91ec", x"91ed", x"91ee", x"91ef", x"91ef", x"91f0", x"91f1", x"91f2", x"91f3",
        x"91f4", x"91f5", x"91f6", x"91f7", x"91f8", x"91f9", x"91f9", x"91fa", x"91fb", x"91fc", x"91fd", x"91fe", x"91ff", x"9200", x"9201", x"9202",
        x"9203", x"9204", x"9205", x"9206", x"9207", x"9208", x"9209", x"920a", x"920b", x"920c", x"920d", x"920e", x"920f", x"9210", x"9211", x"9212",
        x"9213", x"9214", x"9215", x"9216", x"9217", x"9219", x"921a", x"921b", x"921c", x"921d", x"921e", x"921f", x"9220", x"9221", x"9222", x"9224",
        x"9225", x"9226", x"9227", x"9228", x"9229", x"922a", x"922b", x"922d", x"922e", x"922f", x"9230", x"9231", x"9233", x"9234", x"9235", x"9236",
        x"9237", x"9239", x"923a", x"923b", x"923c", x"923d", x"923f", x"9240", x"9241", x"9242", x"9244", x"9245", x"9246", x"9248", x"9249", x"924a",
        x"924b", x"924d", x"924e", x"924f", x"9251", x"9252", x"9253", x"9255", x"9256", x"9257", x"9259", x"925a", x"925b", x"925d", x"925e", x"925f",
        x"9261", x"9262", x"9264", x"9265", x"9266", x"9268", x"9269", x"926b", x"926c", x"926d", x"926f", x"9270", x"9272", x"9273", x"9275", x"9276",
        x"9278", x"9279", x"927a", x"927c", x"927d", x"927f", x"9280", x"9282", x"9283", x"9285", x"9287", x"9288", x"928a", x"928b", x"928d", x"928e",
        x"9290", x"9291", x"9293", x"9294", x"9296", x"9298", x"9299", x"929b", x"929c", x"929e", x"92a0", x"92a1", x"92a3", x"92a5", x"92a6", x"92a8",
        x"92aa", x"92ab", x"92ad", x"92af", x"92b0", x"92b2", x"92b4", x"92b5", x"92b7", x"92b9", x"92ba", x"92bc", x"92be", x"92c0", x"92c1", x"92c3",
        x"92c5", x"92c7", x"92c8", x"92ca", x"92cc", x"92ce", x"92cf", x"92d1", x"92d3", x"92d5", x"92d7", x"92d8", x"92da", x"92dc", x"92de", x"92e0",
        x"92e2", x"92e4", x"92e5", x"92e7", x"92e9", x"92eb", x"92ed", x"92ef", x"92f1", x"92f3", x"92f5", x"92f6", x"92f8", x"92fa", x"92fc", x"92fe",
        x"9300", x"9302", x"9304", x"9306", x"9308", x"930a", x"930c", x"930e", x"9310", x"9312", x"9314", x"9316", x"9318", x"931a", x"931c", x"931e",
        x"9320", x"9322", x"9325", x"9327", x"9329", x"932b", x"932d", x"932f", x"9331", x"9333", x"9335", x"9338", x"933a", x"933c", x"933e", x"9340",
        x"9342", x"9345", x"9347", x"9349", x"934b", x"934d", x"9350", x"9352", x"9354", x"9356", x"9358", x"935b", x"935d", x"935f", x"9362", x"9364",
        x"9366", x"9368", x"936b", x"936d", x"936f", x"9372", x"9374", x"9376", x"9379", x"937b", x"937d", x"9380", x"9382", x"9384", x"9387", x"9389",
        x"938c", x"938e", x"9390", x"9393", x"9395", x"9398", x"939a", x"939d", x"939f", x"93a2", x"93a4", x"93a7", x"93a9", x"93ac", x"93ae", x"93b1",
        x"93b3", x"93b6", x"93b8", x"93bb", x"93bd", x"93c0", x"93c2", x"93c5", x"93c8", x"93ca", x"93cd", x"93cf", x"93d2", x"93d5", x"93d7", x"93da",
        x"93dc", x"93df", x"93e2", x"93e4", x"93e7", x"93ea", x"93ed", x"93ef", x"93f2", x"93f5", x"93f7", x"93fa", x"93fd", x"9400", x"9402", x"9405",
        x"9408", x"940b", x"940d", x"9410", x"9413", x"9416", x"9419", x"941c", x"941e", x"9421", x"9424", x"9427", x"942a", x"942d", x"9430", x"9432",
        x"9435", x"9438", x"943b", x"943e", x"9441", x"9444", x"9447", x"944a", x"944d", x"9450", x"9453", x"9456", x"9459", x"945c", x"945f", x"9462",
        x"9465", x"9468", x"946b", x"946e", x"9471", x"9474", x"9477", x"947a", x"947d", x"9480", x"9484", x"9487", x"948a", x"948d", x"9490", x"9493",
        x"9496", x"949a", x"949d", x"94a0", x"94a3", x"94a6", x"94aa", x"94ad", x"94b0", x"94b3", x"94b7", x"94ba", x"94bd", x"94c0", x"94c4", x"94c7",
        x"94ca", x"94ce", x"94d1", x"94d4", x"94d8", x"94db", x"94de", x"94e2", x"94e5", x"94e8", x"94ec", x"94ef", x"94f3", x"94f6", x"94fa", x"94fd",
        x"9500", x"9504", x"9507", x"950b", x"950e", x"9512", x"9515", x"9519", x"951c", x"9520", x"9523", x"9527", x"952b", x"952e", x"9532", x"9535",
        x"9539", x"953c", x"9540", x"9544", x"9547", x"954b", x"954f", x"9552", x"9556", x"955a", x"955d", x"9561", x"9565", x"9568", x"956c", x"9570",
        x"9574", x"9577", x"957b", x"957f", x"9583", x"9586", x"958a", x"958e", x"9592", x"9596", x"959a", x"959d", x"95a1", x"95a5", x"95a9", x"95ad",
        x"95b1", x"95b5", x"95b9", x"95bc", x"95c0", x"95c4", x"95c8", x"95cc", x"95d0", x"95d4", x"95d8", x"95dc", x"95e0", x"95e4", x"95e8", x"95ec",
        x"95f0", x"95f4", x"95f8", x"95fd", x"9601", x"9605", x"9609", x"960d", x"9611", x"9615", x"9619", x"961d", x"9622", x"9626", x"962a", x"962e",
        x"9632", x"9637", x"963b", x"963f", x"9643", x"9648", x"964c", x"9650", x"9654", x"9659", x"965d", x"9661", x"9666", x"966a", x"966e", x"9673",
        x"9677", x"967b", x"9680", x"9684", x"9689", x"968d", x"9691", x"9696", x"969a", x"969f", x"96a3", x"96a8", x"96ac", x"96b1", x"96b5", x"96ba",
        x"96be", x"96c3", x"96c7", x"96cc", x"96d1", x"96d5", x"96da", x"96de", x"96e3", x"96e8", x"96ec", x"96f1", x"96f5", x"96fa", x"96ff", x"9704",
        x"9708", x"970d", x"9712", x"9716", x"971b", x"9720", x"9725", x"9729", x"972e", x"9733", x"9738", x"973d", x"9741", x"9746", x"974b", x"9750",
        x"9755", x"975a", x"975f", x"9763", x"9768", x"976d", x"9772", x"9777", x"977c", x"9781", x"9786", x"978b", x"9790", x"9795", x"979a", x"979f",
        x"97a4", x"97a9", x"97ae", x"97b3", x"97b8", x"97be", x"97c3", x"97c8", x"97cd", x"97d2", x"97d7", x"97dc", x"97e2", x"97e7", x"97ec", x"97f1",
        x"97f6", x"97fc", x"9801", x"9806", x"980b", x"9811", x"9816", x"981b", x"9820", x"9826", x"982b", x"9830", x"9836", x"983b", x"9841", x"9846",
        x"984b", x"9851", x"9856", x"985c", x"9861", x"9867", x"986c", x"9871", x"9877", x"987c", x"9882", x"9887", x"988d", x"9893", x"9898", x"989e",
        x"98a3", x"98a9", x"98ae", x"98b4", x"98ba", x"98bf", x"98c5", x"98cb", x"98d0", x"98d6", x"98dc", x"98e1", x"98e7", x"98ed", x"98f3", x"98f8",
        x"98fe", x"9904", x"990a", x"990f", x"9915", x"991b", x"9921", x"9927", x"992d", x"9933", x"9938", x"993e", x"9944", x"994a", x"9950", x"9956",
        x"995c", x"9962", x"9968", x"996e", x"9974", x"997a", x"9980", x"9986", x"998c", x"9992", x"9998", x"999e", x"99a4", x"99aa", x"99b1", x"99b7",
        x"99bd", x"99c3", x"99c9", x"99cf", x"99d6", x"99dc", x"99e2", x"99e8", x"99ee", x"99f5", x"99fb", x"9a01", x"9a08", x"9a0e", x"9a14", x"9a1b",
        x"9a21", x"9a27", x"9a2e", x"9a34", x"9a3a", x"9a41", x"9a47", x"9a4e", x"9a54", x"9a5a", x"9a61", x"9a67", x"9a6e", x"9a74", x"9a7b", x"9a81",
        x"9a88", x"9a8f", x"9a95", x"9a9c", x"9aa2", x"9aa9", x"9aaf", x"9ab6", x"9abd", x"9ac3", x"9aca", x"9ad1", x"9ad7", x"9ade", x"9ae5", x"9aec",
        x"9af2", x"9af9", x"9b00", x"9b07", x"9b0d", x"9b14", x"9b1b", x"9b22", x"9b29", x"9b2f", x"9b36", x"9b3d", x"9b44", x"9b4b", x"9b52", x"9b59",
        x"9b60", x"9b67", x"9b6e", x"9b75", x"9b7c", x"9b83", x"9b8a", x"9b91", x"9b98", x"9b9f", x"9ba6", x"9bad", x"9bb4", x"9bbb", x"9bc2", x"9bc9",
        x"9bd1", x"9bd8", x"9bdf", x"9be6", x"9bed", x"9bf5", x"9bfc", x"9c03", x"9c0a", x"9c11", x"9c19", x"9c20", x"9c27", x"9c2f", x"9c36", x"9c3d",
        x"9c45", x"9c4c", x"9c53", x"9c5b", x"9c62", x"9c6a", x"9c71", x"9c79", x"9c80", x"9c87", x"9c8f", x"9c96", x"9c9e", x"9ca5", x"9cad", x"9cb5",
        x"9cbc", x"9cc4", x"9ccb", x"9cd3", x"9cdb", x"9ce2", x"9cea", x"9cf1", x"9cf9", x"9d01", x"9d08", x"9d10", x"9d18", x"9d20", x"9d27", x"9d2f",
        x"9d37", x"9d3f", x"9d47", x"9d4e", x"9d56", x"9d5e", x"9d66", x"9d6e", x"9d76", x"9d7e", x"9d85", x"9d8d", x"9d95", x"9d9d", x"9da5", x"9dad",
        x"9db5", x"9dbd", x"9dc5", x"9dcd", x"9dd5", x"9ddd", x"9de5", x"9dee", x"9df6", x"9dfe", x"9e06", x"9e0e", x"9e16", x"9e1e", x"9e27", x"9e2f",
        x"9e37", x"9e3f", x"9e47", x"9e50", x"9e58", x"9e60", x"9e68", x"9e71", x"9e79", x"9e81", x"9e8a", x"9e92", x"9e9b", x"9ea3", x"9eab", x"9eb4",
        x"9ebc", x"9ec5", x"9ecd", x"9ed6", x"9ede", x"9ee7", x"9eef", x"9ef8", x"9f00", x"9f09", x"9f11", x"9f1a", x"9f22", x"9f2b", x"9f34", x"9f3c",
        x"9f45", x"9f4e", x"9f56", x"9f5f", x"9f68", x"9f70", x"9f79", x"9f82", x"9f8b", x"9f93", x"9f9c", x"9fa5", x"9fae", x"9fb7", x"9fc0", x"9fc8",
        x"9fd1", x"9fda", x"9fe3", x"9fec", x"9ff5", x"9ffe", x"a007", x"a010", x"a019", x"a022", x"a02b", x"a034", x"a03d", x"a046", x"a04f", x"a058",
        x"a061", x"a06a", x"a073", x"a07d", x"a086", x"a08f", x"a098", x"a0a1", x"a0ab", x"a0b4", x"a0bd", x"a0c6", x"a0d0", x"a0d9", x"a0e2", x"a0eb",
        x"a0f5", x"a0fe", x"a107", x"a111", x"a11a", x"a124", x"a12d", x"a136", x"a140", x"a149", x"a153", x"a15c", x"a166", x"a16f", x"a179", x"a182",
        x"a18c", x"a196", x"a19f", x"a1a9", x"a1b2", x"a1bc", x"a1c6", x"a1cf", x"a1d9", x"a1e3", x"a1ec", x"a1f6", x"a200", x"a20a", x"a213", x"a21d",
        x"a227", x"a231", x"a23b", x"a244", x"a24e", x"a258", x"a262", x"a26c", x"a276", x"a280", x"a28a", x"a294", x"a29e", x"a2a8", x"a2b2", x"a2bc",
        x"a2c6", x"a2d0", x"a2da", x"a2e4", x"a2ee", x"a2f8", x"a302", x"a30c", x"a316", x"a321", x"a32b", x"a335", x"a33f", x"a349", x"a354", x"a35e",
        x"a368", x"a372", x"a37d", x"a387", x"a391", x"a39c", x"a3a6", x"a3b0", x"a3bb", x"a3c5", x"a3cf", x"a3da", x"a3e4", x"a3ef", x"a3f9", x"a404",
        x"a40e", x"a419", x"a423", x"a42e", x"a438", x"a443", x"a44e", x"a458", x"a463", x"a46d", x"a478", x"a483", x"a48d", x"a498", x"a4a3", x"a4ae",
        x"a4b8", x"a4c3", x"a4ce", x"a4d9", x"a4e3", x"a4ee", x"a4f9", x"a504", x"a50f", x"a51a", x"a524", x"a52f", x"a53a", x"a545", x"a550", x"a55b",
        x"a566", x"a571", x"a57c", x"a587", x"a592", x"a59d", x"a5a8", x"a5b3", x"a5be", x"a5ca", x"a5d5", x"a5e0", x"a5eb", x"a5f6", x"a601", x"a60d",
        x"a618", x"a623", x"a62e", x"a639", x"a645", x"a650", x"a65b", x"a667", x"a672", x"a67d", x"a689", x"a694", x"a6a0", x"a6ab", x"a6b6", x"a6c2",
        x"a6cd", x"a6d9", x"a6e4", x"a6f0", x"a6fb", x"a707", x"a712", x"a71e", x"a729", x"a735", x"a741", x"a74c", x"a758", x"a764", x"a76f", x"a77b",
        x"a787", x"a792", x"a79e", x"a7aa", x"a7b6", x"a7c1", x"a7cd", x"a7d9", x"a7e5", x"a7f1", x"a7fd", x"a808", x"a814", x"a820", x"a82c", x"a838",
        x"a844", x"a850", x"a85c", x"a868", x"a874", x"a880", x"a88c", x"a898", x"a8a4", x"a8b0", x"a8bc", x"a8c8", x"a8d5", x"a8e1", x"a8ed", x"a8f9",
        x"a905", x"a911", x"a91e", x"a92a", x"a936", x"a942", x"a94f", x"a95b", x"a967", x"a974", x"a980", x"a98c", x"a999", x"a9a5", x"a9b1", x"a9be",
        x"a9ca", x"a9d7", x"a9e3", x"a9f0", x"a9fc", x"aa09", x"aa15", x"aa22", x"aa2e", x"aa3b", x"aa48", x"aa54", x"aa61", x"aa6d", x"aa7a", x"aa87",
        x"aa93", x"aaa0", x"aaad", x"aab9", x"aac6", x"aad3", x"aae0", x"aaed", x"aaf9", x"ab06", x"ab13", x"ab20", x"ab2d", x"ab3a", x"ab47", x"ab53",
        x"ab60", x"ab6d", x"ab7a", x"ab87", x"ab94", x"aba1", x"abae", x"abbb", x"abc8", x"abd5", x"abe2", x"abf0", x"abfd", x"ac0a", x"ac17", x"ac24",
        x"ac31", x"ac3e", x"ac4c", x"ac59", x"ac66", x"ac73", x"ac81", x"ac8e", x"ac9b", x"aca9", x"acb6", x"acc3", x"acd1", x"acde", x"aceb", x"acf9",
        x"ad06", x"ad14", x"ad21", x"ad2f", x"ad3c", x"ad49", x"ad57", x"ad65", x"ad72", x"ad80", x"ad8d", x"ad9b", x"ada8", x"adb6", x"adc4", x"add1",
        x"addf", x"aded", x"adfa", x"ae08", x"ae16", x"ae24", x"ae31", x"ae3f", x"ae4d", x"ae5b", x"ae68", x"ae76", x"ae84", x"ae92", x"aea0", x"aeae",
        x"aebc", x"aeca", x"aed8", x"aee6", x"aef4", x"af02", x"af10", x"af1e", x"af2c", x"af3a", x"af48", x"af56", x"af64", x"af72", x"af80", x"af8e",
        x"af9c", x"afab", x"afb9", x"afc7", x"afd5", x"afe3", x"aff2", x"b000", x"b00e", x"b01d", x"b02b", x"b039", x"b048", x"b056", x"b064", x"b073",
        x"b081", x"b090", x"b09e", x"b0ac", x"b0bb", x"b0c9", x"b0d8", x"b0e6", x"b0f5", x"b103", x"b112", x"b121", x"b12f", x"b13e", x"b14c", x"b15b",
        x"b16a", x"b178", x"b187", x"b196", x"b1a4", x"b1b3", x"b1c2", x"b1d1", x"b1df", x"b1ee", x"b1fd", x"b20c", x"b21b", x"b22a", x"b238", x"b247",
        x"b256", x"b265", x"b274", x"b283", x"b292", x"b2a1", x"b2b0", x"b2bf", x"b2ce", x"b2dd", x"b2ec", x"b2fb", x"b30a", x"b319", x"b328", x"b338",
        x"b347", x"b356", x"b365", x"b374", x"b383", x"b393", x"b3a2", x"b3b1", x"b3c0", x"b3d0", x"b3df", x"b3ee", x"b3fe", x"b40d", x"b41c", x"b42c",
        x"b43b", x"b44a", x"b45a", x"b469", x"b479", x"b488", x"b498", x"b4a7", x"b4b7", x"b4c6", x"b4d6", x"b4e5", x"b4f5", x"b504", x"b514", x"b524",
        x"b533", x"b543", x"b553", x"b562", x"b572", x"b582", x"b591", x"b5a1", x"b5b1", x"b5c1", x"b5d0", x"b5e0", x"b5f0", x"b600", x"b610", x"b620",
        x"b62f", x"b63f", x"b64f", x"b65f", x"b66f", x"b67f", x"b68f", x"b69f", x"b6af", x"b6bf", x"b6cf", x"b6df", x"b6ef", x"b6ff", x"b70f", x"b71f",
        x"b72f", x"b740", x"b750", x"b760", x"b770", x"b780", x"b790", x"b7a1", x"b7b1", x"b7c1", x"b7d1", x"b7e2", x"b7f2", x"b802", x"b813", x"b823",
        x"b833", x"b844", x"b854", x"b864", x"b875", x"b885", x"b896", x"b8a6", x"b8b7", x"b8c7", x"b8d8", x"b8e8", x"b8f9", x"b909", x"b91a", x"b92a",
        x"b93b", x"b94c", x"b95c", x"b96d", x"b97d", x"b98e", x"b99f", x"b9af", x"b9c0", x"b9d1", x"b9e2", x"b9f2", x"ba03", x"ba14", x"ba25", x"ba36",
        x"ba46", x"ba57", x"ba68", x"ba79", x"ba8a", x"ba9b", x"baac", x"babd", x"bacd", x"bade", x"baef", x"bb00", x"bb11", x"bb22", x"bb33", x"bb44",
        x"bb56", x"bb67", x"bb78", x"bb89", x"bb9a", x"bbab", x"bbbc", x"bbcd", x"bbdf", x"bbf0", x"bc01", x"bc12", x"bc23", x"bc35", x"bc46", x"bc57",
        x"bc69", x"bc7a", x"bc8b", x"bc9c", x"bcae", x"bcbf", x"bcd1", x"bce2", x"bcf3", x"bd05", x"bd16", x"bd28", x"bd39", x"bd4b", x"bd5c", x"bd6e",
        x"bd7f", x"bd91", x"bda2", x"bdb4", x"bdc5", x"bdd7", x"bde9", x"bdfa", x"be0c", x"be1e", x"be2f", x"be41", x"be53", x"be64", x"be76", x"be88",
        x"be99", x"beab", x"bebd", x"becf", x"bee1", x"bef2", x"bf04", x"bf16", x"bf28", x"bf3a", x"bf4c", x"bf5e", x"bf70", x"bf82", x"bf94", x"bfa5",
        x"bfb7", x"bfc9", x"bfdb", x"bfed", x"c000", x"c012", x"c024", x"c036", x"c048", x"c05a", x"c06c", x"c07e", x"c090", x"c0a2", x"c0b5", x"c0c7",
        x"c0d9", x"c0eb", x"c0fd", x"c110", x"c122", x"c134", x"c147", x"c159", x"c16b", x"c17d", x"c190", x"c1a2", x"c1b5", x"c1c7", x"c1d9", x"c1ec",
        x"c1fe", x"c211", x"c223", x"c236", x"c248", x"c25a", x"c26d", x"c280", x"c292", x"c2a5", x"c2b7", x"c2ca", x"c2dc", x"c2ef", x"c302", x"c314",
        x"c327", x"c339", x"c34c", x"c35f", x"c372", x"c384", x"c397", x"c3aa", x"c3bc", x"c3cf", x"c3e2", x"c3f5", x"c408", x"c41a", x"c42d", x"c440",
        x"c453", x"c466", x"c479", x"c48c", x"c49f", x"c4b1", x"c4c4", x"c4d7", x"c4ea", x"c4fd", x"c510", x"c523", x"c536", x"c549", x"c55c", x"c56f",
        x"c582", x"c596", x"c5a9", x"c5bc", x"c5cf", x"c5e2", x"c5f5", x"c608", x"c61c", x"c62f", x"c642", x"c655", x"c668", x"c67c", x"c68f", x"c6a2",
        x"c6b5", x"c6c9", x"c6dc", x"c6ef", x"c703", x"c716", x"c729", x"c73d", x"c750", x"c764", x"c777", x"c78a", x"c79e", x"c7b1", x"c7c5", x"c7d8",
        x"c7ec", x"c7ff", x"c813", x"c826", x"c83a", x"c84d", x"c861", x"c875", x"c888", x"c89c", x"c8af", x"c8c3", x"c8d7", x"c8ea", x"c8fe", x"c912",
        x"c925", x"c939", x"c94d", x"c960", x"c974", x"c988", x"c99c", x"c9b0", x"c9c3", x"c9d7", x"c9eb", x"c9ff", x"ca13", x"ca26", x"ca3a", x"ca4e",
        x"ca62", x"ca76", x"ca8a", x"ca9e", x"cab2", x"cac6", x"cada", x"caee", x"cb02", x"cb16", x"cb2a", x"cb3e", x"cb52", x"cb66", x"cb7a", x"cb8e",
        x"cba2", x"cbb6", x"cbca", x"cbde", x"cbf3", x"cc07", x"cc1b", x"cc2f", x"cc43", x"cc57", x"cc6c", x"cc80", x"cc94", x"cca8", x"ccbd", x"ccd1",
        x"cce5", x"ccf9", x"cd0e", x"cd22", x"cd36", x"cd4b", x"cd5f", x"cd74", x"cd88", x"cd9c", x"cdb1", x"cdc5", x"cdda", x"cdee", x"ce02", x"ce17",
        x"ce2b", x"ce40", x"ce54", x"ce69", x"ce7d", x"ce92", x"cea6", x"cebb", x"ced0", x"cee4", x"cef9", x"cf0d", x"cf22", x"cf37", x"cf4b", x"cf60",
        x"cf74", x"cf89", x"cf9e", x"cfb3", x"cfc7", x"cfdc", x"cff1", x"d005", x"d01a", x"d02f", x"d044", x"d058", x"d06d", x"d082", x"d097", x"d0ac",
        x"d0c1", x"d0d5", x"d0ea", x"d0ff", x"d114", x"d129", x"d13e", x"d153", x"d168", x"d17d", x"d192", x"d1a7", x"d1bc", x"d1d1", x"d1e6", x"d1fb",
        x"d210", x"d225", x"d23a", x"d24f", x"d264", x"d279", x"d28e", x"d2a3", x"d2b8", x"d2cd", x"d2e2", x"d2f7", x"d30d", x"d322", x"d337", x"d34c",
        x"d361", x"d377", x"d38c", x"d3a1", x"d3b6", x"d3cb", x"d3e1", x"d3f6", x"d40b", x"d420", x"d436", x"d44b", x"d460", x"d476", x"d48b", x"d4a0",
        x"d4b6", x"d4cb", x"d4e1", x"d4f6", x"d50b", x"d521", x"d536", x"d54c", x"d561", x"d577", x"d58c", x"d5a1", x"d5b7", x"d5cc", x"d5e2", x"d5f7",
        x"d60d", x"d622", x"d638", x"d64e", x"d663", x"d679", x"d68e", x"d6a4", x"d6ba", x"d6cf", x"d6e5", x"d6fa", x"d710", x"d726", x"d73b", x"d751",
        x"d767", x"d77c", x"d792", x"d7a8", x"d7be", x"d7d3", x"d7e9", x"d7ff", x"d815", x"d82a", x"d840", x"d856", x"d86c", x"d881", x"d897", x"d8ad",
        x"d8c3", x"d8d9", x"d8ef", x"d905", x"d91a", x"d930", x"d946", x"d95c", x"d972", x"d988", x"d99e", x"d9b4", x"d9ca", x"d9e0", x"d9f6", x"da0c",
        x"da22", x"da38", x"da4e", x"da64", x"da7a", x"da90", x"daa6", x"dabc", x"dad2", x"dae8", x"dafe", x"db14", x"db2a", x"db40", x"db57", x"db6d",
        x"db83", x"db99", x"dbaf", x"dbc5", x"dbdb", x"dbf2", x"dc08", x"dc1e", x"dc34", x"dc4a", x"dc61", x"dc77", x"dc8d", x"dca3", x"dcba", x"dcd0",
        x"dce6", x"dcfc", x"dd13", x"dd29", x"dd3f", x"dd56", x"dd6c", x"dd82", x"dd99", x"ddaf", x"ddc5", x"dddc", x"ddf2", x"de09", x"de1f", x"de35",
        x"de4c", x"de62", x"de79", x"de8f", x"dea5", x"debc", x"ded2", x"dee9", x"deff", x"df16", x"df2c", x"df43", x"df59", x"df70", x"df86", x"df9d",
        x"dfb3", x"dfca", x"dfe1", x"dff7", x"e00e", x"e024", x"e03b", x"e051", x"e068", x"e07f", x"e095", x"e0ac", x"e0c3", x"e0d9", x"e0f0", x"e107",
        x"e11d", x"e134", x"e14b", x"e161", x"e178", x"e18f", x"e1a5", x"e1bc", x"e1d3", x"e1ea", x"e200", x"e217", x"e22e", x"e245", x"e25b", x"e272",
        x"e289", x"e2a0", x"e2b7", x"e2cd", x"e2e4", x"e2fb", x"e312", x"e329", x"e340", x"e356", x"e36d", x"e384", x"e39b", x"e3b2", x"e3c9", x"e3e0",
        x"e3f7", x"e40d", x"e424", x"e43b", x"e452", x"e469", x"e480", x"e497", x"e4ae", x"e4c5", x"e4dc", x"e4f3", x"e50a", x"e521", x"e538", x"e54f",
        x"e566", x"e57d", x"e594", x"e5ab", x"e5c2", x"e5d9", x"e5f0", x"e607", x"e61e", x"e635", x"e64c", x"e664", x"e67b", x"e692", x"e6a9", x"e6c0",
        x"e6d7", x"e6ee", x"e705", x"e71c", x"e734", x"e74b", x"e762", x"e779", x"e790", x"e7a7", x"e7bf", x"e7d6", x"e7ed", x"e804", x"e81b", x"e833",
        x"e84a", x"e861", x"e878", x"e88f", x"e8a7", x"e8be", x"e8d5", x"e8ec", x"e904", x"e91b", x"e932", x"e949", x"e961", x"e978", x"e98f", x"e9a7",
        x"e9be", x"e9d5", x"e9ed", x"ea04", x"ea1b", x"ea33", x"ea4a", x"ea61", x"ea79", x"ea90", x"eaa7", x"eabf", x"ead6", x"eaed", x"eb05", x"eb1c",
        x"eb34", x"eb4b", x"eb62", x"eb7a", x"eb91", x"eba9", x"ebc0", x"ebd8", x"ebef", x"ec06", x"ec1e", x"ec35", x"ec4d", x"ec64", x"ec7c", x"ec93",
        x"ecab", x"ecc2", x"ecda", x"ecf1", x"ed09", x"ed20", x"ed38", x"ed4f", x"ed67", x"ed7e", x"ed96", x"edad", x"edc5", x"eddc", x"edf4", x"ee0b",
        x"ee23", x"ee3a", x"ee52", x"ee6a", x"ee81", x"ee99", x"eeb0", x"eec8", x"eee0", x"eef7", x"ef0f", x"ef26", x"ef3e", x"ef56", x"ef6d", x"ef85",
        x"ef9c", x"efb4", x"efcc", x"efe3", x"effb", x"f013", x"f02a", x"f042", x"f059", x"f071", x"f089", x"f0a0", x"f0b8", x"f0d0", x"f0e7", x"f0ff",
        x"f117", x"f12f", x"f146", x"f15e", x"f176", x"f18d", x"f1a5", x"f1bd", x"f1d4", x"f1ec", x"f204", x"f21c", x"f233", x"f24b", x"f263", x"f27b",
        x"f292", x"f2aa", x"f2c2", x"f2da", x"f2f1", x"f309", x"f321", x"f339", x"f350", x"f368", x"f380", x"f398", x"f3af", x"f3c7", x"f3df", x"f3f7",
        x"f40f", x"f426", x"f43e", x"f456", x"f46e", x"f486", x"f49d", x"f4b5", x"f4cd", x"f4e5", x"f4fd", x"f515", x"f52c", x"f544", x"f55c", x"f574",
        x"f58c", x"f5a4", x"f5bb", x"f5d3", x"f5eb", x"f603", x"f61b", x"f633", x"f64b", x"f662", x"f67a", x"f692", x"f6aa", x"f6c2", x"f6da", x"f6f2",
        x"f70a", x"f721", x"f739", x"f751", x"f769", x"f781", x"f799", x"f7b1", x"f7c9", x"f7e1", x"f7f8", x"f810", x"f828", x"f840", x"f858", x"f870",
        x"f888", x"f8a0", x"f8b8", x"f8d0", x"f8e8", x"f900", x"f917", x"f92f", x"f947", x"f95f", x"f977", x"f98f", x"f9a7", x"f9bf", x"f9d7", x"f9ef",
        x"fa07", x"fa1f", x"fa37", x"fa4f", x"fa67", x"fa7f", x"fa96", x"faae", x"fac6", x"fade", x"faf6", x"fb0e", x"fb26", x"fb3e", x"fb56", x"fb6e",
        x"fb86", x"fb9e", x"fbb6", x"fbce", x"fbe6", x"fbfe", x"fc16", x"fc2e", x"fc46", x"fc5e", x"fc76", x"fc8e", x"fca6", x"fcbe", x"fcd6", x"fcee",
        x"fd06", x"fd1e", x"fd36", x"fd4e", x"fd66", x"fd7e", x"fd96", x"fdad", x"fdc5", x"fddd", x"fdf5", x"fe0d", x"fe25", x"fe3d", x"fe55", x"fe6d",
        x"fe85", x"fe9d", x"feb5", x"fecd", x"fee5", x"fefd", x"ff15", x"ff2d", x"ff45", x"ff5d", x"ff75", x"ff8d", x"ffa5", x"ffbd", x"ffd5", x"ffed",
        x"0004", x"001c", x"0034", x"004c", x"0064", x"007c", x"0094", x"00ac", x"00c4", x"00dc", x"00f4", x"010c", x"0124", x"013c", x"0154", x"016c",
        x"0184", x"019c", x"01b4", x"01cc", x"01e4", x"01fc", x"0214", x"022c", x"0244", x"025c", x"0274", x"028c", x"02a4", x"02bc", x"02d4", x"02ec",
        x"0304", x"031c", x"0334", x"034c", x"0364", x"037c", x"0394", x"03ac", x"03c4", x"03dc", x"03f4", x"040c", x"0423", x"043b", x"0453", x"046b",
        x"0483", x"049b", x"04b3", x"04cb", x"04e3", x"04fb", x"0513", x"052b", x"0543", x"055b", x"0573", x"058b", x"05a3", x"05bb", x"05d3", x"05eb",
        x"0603", x"061b", x"0632", x"064a", x"0662", x"067a", x"0692", x"06aa", x"06c2", x"06da", x"06f2", x"070a", x"0722", x"073a", x"0752", x"076a",
        x"0781", x"0799", x"07b1", x"07c9", x"07e1", x"07f9", x"0811", x"0829", x"0841", x"0859", x"0870", x"0888", x"08a0", x"08b8", x"08d0", x"08e8",
        x"0900", x"0918", x"0930", x"0947", x"095f", x"0977", x"098f", x"09a7", x"09bf", x"09d7", x"09ef", x"0a06", x"0a1e", x"0a36", x"0a4e", x"0a66",
        x"0a7e", x"0a95", x"0aad", x"0ac5", x"0add", x"0af5", x"0b0d", x"0b24", x"0b3c", x"0b54", x"0b6c", x"0b84", x"0b9b", x"0bb3", x"0bcb", x"0be3",
        x"0bfb", x"0c12", x"0c2a", x"0c42", x"0c5a", x"0c72", x"0c89", x"0ca1", x"0cb9", x"0cd1", x"0ce8", x"0d00", x"0d18", x"0d30", x"0d48", x"0d5f",
        x"0d77", x"0d8f", x"0da6", x"0dbe", x"0dd6", x"0dee", x"0e05", x"0e1d", x"0e35", x"0e4d", x"0e64", x"0e7c", x"0e94", x"0eab", x"0ec3", x"0edb",
        x"0ef2", x"0f0a", x"0f22", x"0f39", x"0f51", x"0f69", x"0f80", x"0f98", x"0fb0", x"0fc7", x"0fdf", x"0ff7", x"100e", x"1026", x"103e", x"1055",
        x"106d", x"1085", x"109c", x"10b4", x"10cb", x"10e3", x"10fb", x"1112", x"112a", x"1141", x"1159", x"1170", x"1188", x"11a0", x"11b7", x"11cf",
        x"11e6", x"11fe", x"1215", x"122d", x"1244", x"125c", x"1274", x"128b", x"12a3", x"12ba", x"12d2", x"12e9", x"1301", x"1318", x"1330", x"1347",
        x"135f", x"1376", x"138d", x"13a5", x"13bc", x"13d4", x"13eb", x"1403", x"141a", x"1432", x"1449", x"1460", x"1478", x"148f", x"14a7", x"14be",
        x"14d6", x"14ed", x"1504", x"151c", x"1533", x"154a", x"1562", x"1579", x"1590", x"15a8", x"15bf", x"15d7", x"15ee", x"1605", x"161d", x"1634",
        x"164b", x"1662", x"167a", x"1691", x"16a8", x"16c0", x"16d7", x"16ee", x"1705", x"171d", x"1734", x"174b", x"1762", x"177a", x"1791", x"17a8",
        x"17bf", x"17d7", x"17ee", x"1805", x"181c", x"1833", x"184b", x"1862", x"1879", x"1890", x"18a7", x"18be", x"18d5", x"18ed", x"1904", x"191b",
        x"1932", x"1949", x"1960", x"1977", x"198e", x"19a5", x"19bd", x"19d4", x"19eb", x"1a02", x"1a19", x"1a30", x"1a47", x"1a5e", x"1a75", x"1a8c",
        x"1aa3", x"1aba", x"1ad1", x"1ae8", x"1aff", x"1b16", x"1b2d", x"1b44", x"1b5b", x"1b72", x"1b89", x"1ba0", x"1bb7", x"1bce", x"1be5", x"1bfb",
        x"1c12", x"1c29", x"1c40", x"1c57", x"1c6e", x"1c85", x"1c9c", x"1cb3", x"1cc9", x"1ce0", x"1cf7", x"1d0e", x"1d25", x"1d3c", x"1d52", x"1d69",
        x"1d80", x"1d97", x"1dad", x"1dc4", x"1ddb", x"1df2", x"1e09", x"1e1f", x"1e36", x"1e4d", x"1e63", x"1e7a", x"1e91", x"1ea8", x"1ebe", x"1ed5",
        x"1eec", x"1f02", x"1f19", x"1f30", x"1f46", x"1f5d", x"1f73", x"1f8a", x"1fa1", x"1fb7", x"1fce", x"1fe4", x"1ffb", x"2012", x"2028", x"203f",
        x"2055", x"206c", x"2082", x"2099", x"20af", x"20c6", x"20dc", x"20f3", x"2109", x"2120", x"2136", x"214d", x"2163", x"217a", x"2190", x"21a7",
        x"21bd", x"21d3", x"21ea", x"2200", x"2217", x"222d", x"2243", x"225a", x"2270", x"2286", x"229d", x"22b3", x"22c9", x"22e0", x"22f6", x"230c",
        x"2322", x"2339", x"234f", x"2365", x"237b", x"2392", x"23a8", x"23be", x"23d4", x"23eb", x"2401", x"2417", x"242d", x"2443", x"2459", x"2470",
        x"2486", x"249c", x"24b2", x"24c8", x"24de", x"24f4", x"250a", x"2520", x"2537", x"254d", x"2563", x"2579", x"258f", x"25a5", x"25bb", x"25d1",
        x"25e7", x"25fd", x"2613", x"2629", x"263f", x"2655", x"266b", x"2680", x"2696", x"26ac", x"26c2", x"26d8", x"26ee", x"2704", x"271a", x"2730",
        x"2745", x"275b", x"2771", x"2787", x"279d", x"27b3", x"27c8", x"27de", x"27f4", x"280a", x"281f", x"2835", x"284b", x"2861", x"2876", x"288c",
        x"28a2", x"28b7", x"28cd", x"28e3", x"28f8", x"290e", x"2924", x"2939", x"294f", x"2964", x"297a", x"2990", x"29a5", x"29bb", x"29d0", x"29e6",
        x"29fb", x"2a11", x"2a26", x"2a3c", x"2a51", x"2a67", x"2a7c", x"2a92", x"2aa7", x"2abd", x"2ad2", x"2ae7", x"2afd", x"2b12", x"2b28", x"2b3d",
        x"2b52", x"2b68", x"2b7d", x"2b92", x"2ba8", x"2bbd", x"2bd2", x"2be8", x"2bfd", x"2c12", x"2c27", x"2c3d", x"2c52", x"2c67", x"2c7c", x"2c92",
        x"2ca7", x"2cbc", x"2cd1", x"2ce6", x"2cfb", x"2d11", x"2d26", x"2d3b", x"2d50", x"2d65", x"2d7a", x"2d8f", x"2da4", x"2db9", x"2dce", x"2de3",
        x"2df8", x"2e0d", x"2e22", x"2e37", x"2e4c", x"2e61", x"2e76", x"2e8b", x"2ea0", x"2eb5", x"2eca", x"2edf", x"2ef4", x"2f09", x"2f1e", x"2f33",
        x"2f47", x"2f5c", x"2f71", x"2f86", x"2f9b", x"2faf", x"2fc4", x"2fd9", x"2fee", x"3002", x"3017", x"302c", x"3041", x"3055", x"306a", x"307f",
        x"3093", x"30a8", x"30bd", x"30d1", x"30e6", x"30fb", x"310f", x"3124", x"3138", x"314d", x"3161", x"3176", x"318a", x"319f", x"31b3", x"31c8",
        x"31dc", x"31f1", x"3205", x"321a", x"322e", x"3243", x"3257", x"326b", x"3280", x"3294", x"32a9", x"32bd", x"32d1", x"32e6", x"32fa", x"330e",
        x"3322", x"3337", x"334b", x"335f", x"3374", x"3388", x"339c", x"33b0", x"33c4", x"33d9", x"33ed", x"3401", x"3415", x"3429", x"343d", x"3451",
        x"3466", x"347a", x"348e", x"34a2", x"34b6", x"34ca", x"34de", x"34f2", x"3506", x"351a", x"352e", x"3542", x"3556", x"356a", x"357e", x"3591",
        x"35a5", x"35b9", x"35cd", x"35e1", x"35f5", x"3609", x"361d", x"3630", x"3644", x"3658", x"366c", x"367f", x"3693", x"36a7", x"36bb", x"36ce",
        x"36e2", x"36f6", x"3709", x"371d", x"3731", x"3744", x"3758", x"376c", x"377f", x"3793", x"37a6", x"37ba", x"37ce", x"37e1", x"37f5", x"3808",
        x"381c", x"382f", x"3843", x"3856", x"3869", x"387d", x"3890", x"38a4", x"38b7", x"38ca", x"38de", x"38f1", x"3905", x"3918", x"392b", x"393e",
        x"3952", x"3965", x"3978", x"398c", x"399f", x"39b2", x"39c5", x"39d8", x"39ec", x"39ff", x"3a12", x"3a25", x"3a38", x"3a4b", x"3a5e", x"3a72",
        x"3a85", x"3a98", x"3aab", x"3abe", x"3ad1", x"3ae4", x"3af7", x"3b0a", x"3b1d", x"3b30", x"3b43", x"3b56", x"3b69", x"3b7b", x"3b8e", x"3ba1",
        x"3bb4", x"3bc7", x"3bda", x"3bed", x"3bff", x"3c12", x"3c25", x"3c38", x"3c4b", x"3c5d", x"3c70", x"3c83", x"3c95", x"3ca8", x"3cbb", x"3ccd",
        x"3ce0", x"3cf3", x"3d05", x"3d18", x"3d2b", x"3d3d", x"3d50", x"3d62", x"3d75", x"3d87", x"3d9a", x"3dac", x"3dbf", x"3dd1", x"3de4", x"3df6",
        x"3e09", x"3e1b", x"3e2d", x"3e40", x"3e52", x"3e65", x"3e77", x"3e89", x"3e9c", x"3eae", x"3ec0", x"3ed3", x"3ee5", x"3ef7", x"3f09", x"3f1b",
        x"3f2e", x"3f40", x"3f52", x"3f64", x"3f76", x"3f89", x"3f9b", x"3fad", x"3fbf", x"3fd1", x"3fe3", x"3ff5", x"4007", x"4019", x"402b", x"403d",
        x"404f", x"4061", x"4073", x"4085", x"4097", x"40a9", x"40bb", x"40cd", x"40df", x"40f0", x"4102", x"4114", x"4126", x"4138", x"4149", x"415b",
        x"416d", x"417f", x"4191", x"41a2", x"41b4", x"41c6", x"41d7", x"41e9", x"41fb", x"420c", x"421e", x"422f", x"4241", x"4253", x"4264", x"4276",
        x"4287", x"4299", x"42aa", x"42bc", x"42cd", x"42df", x"42f0", x"4302", x"4313", x"4324", x"4336", x"4347", x"4359", x"436a", x"437b", x"438c",
        x"439e", x"43af", x"43c0", x"43d2", x"43e3", x"43f4", x"4405", x"4416", x"4428", x"4439", x"444a", x"445b", x"446c", x"447d", x"448e", x"44a0",
        x"44b1", x"44c2", x"44d3", x"44e4", x"44f5", x"4506", x"4517", x"4528", x"4539", x"454a", x"455b", x"456b", x"457c", x"458d", x"459e", x"45af",
        x"45c0", x"45d1", x"45e1", x"45f2", x"4603", x"4614", x"4624", x"4635", x"4646", x"4657", x"4667", x"4678", x"4689", x"4699", x"46aa", x"46ba",
        x"46cb", x"46dc", x"46ec", x"46fd", x"470d", x"471e", x"472e", x"473f", x"474f", x"4760", x"4770", x"4781", x"4791", x"47a1", x"47b2", x"47c2",
        x"47d3", x"47e3", x"47f3", x"4804", x"4814", x"4824", x"4834", x"4845", x"4855", x"4865", x"4875", x"4886", x"4896", x"48a6", x"48b6", x"48c6",
        x"48d6", x"48e6", x"48f7", x"4907", x"4917", x"4927", x"4937", x"4947", x"4957", x"4967", x"4977", x"4987", x"4997", x"49a7", x"49b6", x"49c6",
        x"49d6", x"49e6", x"49f6", x"4a06", x"4a16", x"4a25", x"4a35", x"4a45", x"4a55", x"4a64", x"4a74", x"4a84", x"4a94", x"4aa3", x"4ab3", x"4ac3",
        x"4ad2", x"4ae2", x"4af1", x"4b01", x"4b11", x"4b20", x"4b30", x"4b3f", x"4b4f", x"4b5e", x"4b6e", x"4b7d", x"4b8d", x"4b9c", x"4bac", x"4bbb",
        x"4bca", x"4bda", x"4be9", x"4bf8", x"4c08", x"4c17", x"4c26", x"4c36", x"4c45", x"4c54", x"4c63", x"4c73", x"4c82", x"4c91", x"4ca0", x"4caf",
        x"4cbf", x"4cce", x"4cdd", x"4cec", x"4cfb", x"4d0a", x"4d19", x"4d28", x"4d37", x"4d46", x"4d55", x"4d64", x"4d73", x"4d82", x"4d91", x"4da0",
        x"4daf", x"4dbe", x"4dcd", x"4ddc", x"4dea", x"4df9", x"4e08", x"4e17", x"4e26", x"4e34", x"4e43", x"4e52", x"4e61", x"4e6f", x"4e7e", x"4e8d",
        x"4e9b", x"4eaa", x"4eb9", x"4ec7", x"4ed6", x"4ee4", x"4ef3", x"4f02", x"4f10", x"4f1f", x"4f2d", x"4f3c", x"4f4a", x"4f59", x"4f67", x"4f75",
        x"4f84", x"4f92", x"4fa1", x"4faf", x"4fbd", x"4fcc", x"4fda", x"4fe8", x"4ff7", x"5005", x"5013", x"5021", x"5030", x"503e", x"504c", x"505a",
        x"5068", x"5077", x"5085", x"5093", x"50a1", x"50af", x"50bd", x"50cb", x"50d9", x"50e7", x"50f5", x"5103", x"5111", x"511f", x"512d", x"513b",
        x"5149", x"5157", x"5165", x"5173", x"5181", x"518e", x"519c", x"51aa", x"51b8", x"51c6", x"51d3", x"51e1", x"51ef", x"51fd", x"520a", x"5218",
        x"5226", x"5233", x"5241", x"524f", x"525c", x"526a", x"5277", x"5285", x"5293", x"52a0", x"52ae", x"52bb", x"52c9", x"52d6", x"52e4", x"52f1",
        x"52fe", x"530c", x"5319", x"5327", x"5334", x"5341", x"534f", x"535c", x"5369", x"5377", x"5384", x"5391", x"539e", x"53ac", x"53b9", x"53c6",
        x"53d3", x"53e0", x"53ed", x"53fb", x"5408", x"5415", x"5422", x"542f", x"543c", x"5449", x"5456", x"5463", x"5470", x"547d", x"548a", x"5497",
        x"54a4", x"54b1", x"54be", x"54cb", x"54d8", x"54e4", x"54f1", x"54fe", x"550b", x"5518", x"5524", x"5531", x"553e", x"554b", x"5557", x"5564",
        x"5571", x"557e", x"558a", x"5597", x"55a3", x"55b0", x"55bd", x"55c9", x"55d6", x"55e2", x"55ef", x"55fb", x"5608", x"5614", x"5621", x"562d",
        x"563a", x"5646", x"5653", x"565f", x"566b", x"5678", x"5684", x"5690", x"569d", x"56a9", x"56b5", x"56c2", x"56ce", x"56da", x"56e6", x"56f3",
        x"56ff", x"570b", x"5717", x"5723", x"572f", x"573c", x"5748", x"5754", x"5760", x"576c", x"5778", x"5784", x"5790", x"579c", x"57a8", x"57b4",
        x"57c0", x"57cc", x"57d8", x"57e4", x"57f0", x"57fb", x"5807", x"5813", x"581f", x"582b", x"5837", x"5842", x"584e", x"585a", x"5866", x"5871",
        x"587d", x"5889", x"5894", x"58a0", x"58ac", x"58b7", x"58c3", x"58cf", x"58da", x"58e6", x"58f1", x"58fd", x"5908", x"5914", x"591f", x"592b",
        x"5936", x"5942", x"594d", x"5959", x"5964", x"5970", x"597b", x"5986", x"5992", x"599d", x"59a8", x"59b4", x"59bf", x"59ca", x"59d5", x"59e1",
        x"59ec", x"59f7", x"5a02", x"5a0d", x"5a19", x"5a24", x"5a2f", x"5a3a", x"5a45", x"5a50", x"5a5b", x"5a66", x"5a71", x"5a7c", x"5a87", x"5a92",
        x"5a9d", x"5aa8", x"5ab3", x"5abe", x"5ac9", x"5ad4", x"5adf", x"5aea", x"5af5", x"5b00", x"5b0a", x"5b15", x"5b20", x"5b2b", x"5b36", x"5b40",
        x"5b4b", x"5b56", x"5b61", x"5b6b", x"5b76", x"5b81", x"5b8b", x"5b96", x"5ba1", x"5bab", x"5bb6", x"5bc0", x"5bcb", x"5bd5", x"5be0", x"5bea",
        x"5bf5", x"5bff", x"5c0a", x"5c14", x"5c1f", x"5c29", x"5c34", x"5c3e", x"5c49", x"5c53", x"5c5d", x"5c68", x"5c72", x"5c7c", x"5c87", x"5c91",
        x"5c9b", x"5ca5", x"5cb0", x"5cba", x"5cc4", x"5cce", x"5cd8", x"5ce3", x"5ced", x"5cf7", x"5d01", x"5d0b", x"5d15", x"5d1f", x"5d29", x"5d33",
        x"5d3d", x"5d47", x"5d51", x"5d5b", x"5d65", x"5d6f", x"5d79", x"5d83", x"5d8d", x"5d97", x"5da1", x"5dab", x"5db5", x"5dbf", x"5dc8", x"5dd2",
        x"5ddc", x"5de6", x"5df0", x"5df9", x"5e03", x"5e0d", x"5e16", x"5e20", x"5e2a", x"5e34", x"5e3d", x"5e47", x"5e50", x"5e5a", x"5e64", x"5e6d",
        x"5e77", x"5e80", x"5e8a", x"5e93", x"5e9d", x"5ea6", x"5eb0", x"5eb9", x"5ec3", x"5ecc", x"5ed6", x"5edf", x"5ee9", x"5ef2", x"5efb", x"5f05",
        x"5f0e", x"5f17", x"5f21", x"5f2a", x"5f33", x"5f3c", x"5f46", x"5f4f", x"5f58", x"5f61", x"5f6b", x"5f74", x"5f7d", x"5f86", x"5f8f", x"5f98",
        x"5fa1", x"5fab", x"5fb4", x"5fbd", x"5fc6", x"5fcf", x"5fd8", x"5fe1", x"5fea", x"5ff3", x"5ffc", x"6005", x"600e", x"6017", x"6020", x"6028",
        x"6031", x"603a", x"6043", x"604c", x"6055", x"605e", x"6066", x"606f", x"6078", x"6081", x"6089", x"6092", x"609b", x"60a4", x"60ac", x"60b5",
        x"60be", x"60c6", x"60cf", x"60d7", x"60e0", x"60e9", x"60f1", x"60fa", x"6102", x"610b", x"6113", x"611c", x"6124", x"612d", x"6135", x"613e",
        x"6146", x"614f", x"6157", x"615f", x"6168", x"6170", x"6179", x"6181", x"6189", x"6192", x"619a", x"61a2", x"61aa", x"61b3", x"61bb", x"61c3",
        x"61cb", x"61d4", x"61dc", x"61e4", x"61ec", x"61f4", x"61fc", x"6204", x"620d", x"6215", x"621d", x"6225", x"622d", x"6235", x"623d", x"6245",
        x"624d", x"6255", x"625d", x"6265", x"626d", x"6275", x"627d", x"6285", x"628c", x"6294", x"629c", x"62a4", x"62ac", x"62b4", x"62bc", x"62c3",
        x"62cb", x"62d3", x"62db", x"62e2", x"62ea", x"62f2", x"62fa", x"6301", x"6309", x"6311", x"6318", x"6320", x"6328", x"632f", x"6337", x"633e",
        x"6346", x"634d", x"6355", x"635d", x"6364", x"636c", x"6373", x"637b", x"6382", x"6389", x"6391", x"6398", x"63a0", x"63a7", x"63ae", x"63b6",
        x"63bd", x"63c5", x"63cc", x"63d3", x"63db", x"63e2", x"63e9", x"63f0", x"63f8", x"63ff", x"6406", x"640d", x"6415", x"641c", x"6423", x"642a",
        x"6431", x"6438", x"643f", x"6447", x"644e", x"6455", x"645c", x"6463", x"646a", x"6471", x"6478", x"647f", x"6486", x"648d", x"6494", x"649b",
        x"64a2", x"64a9", x"64b0", x"64b7", x"64be", x"64c4", x"64cb", x"64d2", x"64d9", x"64e0", x"64e7", x"64ee", x"64f4", x"64fb", x"6502", x"6509",
        x"650f", x"6516", x"651d", x"6524", x"652a", x"6531", x"6538", x"653e", x"6545", x"654c", x"6552", x"6559", x"655f", x"6566", x"656c", x"6573",
        x"657a", x"6580", x"6587", x"658d", x"6594", x"659a", x"65a1", x"65a7", x"65ad", x"65b4", x"65ba", x"65c1", x"65c7", x"65ce", x"65d4", x"65da",
        x"65e1", x"65e7", x"65ed", x"65f4", x"65fa", x"6600", x"6606", x"660d", x"6613", x"6619", x"661f", x"6626", x"662c", x"6632", x"6638", x"663e",
        x"6645", x"664b", x"6651", x"6657", x"665d", x"6663", x"6669", x"666f", x"6675", x"667b", x"6681", x"6687", x"668d", x"6693", x"6699", x"669f",
        x"66a5", x"66ab", x"66b1", x"66b7", x"66bd", x"66c3", x"66c9", x"66cf", x"66d5", x"66da", x"66e0", x"66e6", x"66ec", x"66f2", x"66f8", x"66fd",
        x"6703", x"6709", x"670f", x"6714", x"671a", x"6720", x"6726", x"672b", x"6731", x"6737", x"673c", x"6742", x"6747", x"674d", x"6753", x"6758",
        x"675e", x"6763", x"6769", x"676f", x"6774", x"677a", x"677f", x"6785", x"678a", x"6790", x"6795", x"679b", x"67a0", x"67a6", x"67ab", x"67b0",
        x"67b6", x"67bb", x"67c1", x"67c6", x"67cb", x"67d1", x"67d6", x"67db", x"67e1", x"67e6", x"67eb", x"67f0", x"67f6", x"67fb", x"6800", x"6805",
        x"680b", x"6810", x"6815", x"681a", x"681f", x"6825", x"682a", x"682f", x"6834", x"6839", x"683e", x"6843", x"6849", x"684e", x"6853", x"6858",
        x"685d", x"6862", x"6867", x"686c", x"6871", x"6876", x"687b", x"6880", x"6885", x"688a", x"688f", x"6894", x"6899", x"689d", x"68a2", x"68a7",
        x"68ac", x"68b1", x"68b6", x"68bb", x"68bf", x"68c4", x"68c9", x"68ce", x"68d3", x"68d7", x"68dc", x"68e1", x"68e6", x"68ea", x"68ef", x"68f4",
        x"68f9", x"68fd", x"6902", x"6907", x"690b", x"6910", x"6915", x"6919", x"691e", x"6922", x"6927", x"692c", x"6930", x"6935", x"6939", x"693e",
        x"6942", x"6947", x"694c", x"6950", x"6955", x"6959", x"695d", x"6962", x"6966", x"696b", x"696f", x"6974", x"6978", x"697d", x"6981", x"6985",
        x"698a", x"698e", x"6992", x"6997", x"699b", x"699f", x"69a4", x"69a8", x"69ac", x"69b1", x"69b5", x"69b9", x"69bd", x"69c2", x"69c6", x"69ca",
        x"69ce", x"69d2", x"69d7", x"69db", x"69df", x"69e3", x"69e7", x"69eb", x"69f0", x"69f4", x"69f8", x"69fc", x"6a00", x"6a04", x"6a08", x"6a0c",
        x"6a10", x"6a14", x"6a18", x"6a1c", x"6a20", x"6a24", x"6a28", x"6a2c", x"6a30", x"6a34", x"6a38", x"6a3c", x"6a40", x"6a44", x"6a48", x"6a4c",
        x"6a50", x"6a54", x"6a58", x"6a5b", x"6a5f", x"6a63", x"6a67", x"6a6b", x"6a6f", x"6a72", x"6a76", x"6a7a", x"6a7e", x"6a82", x"6a85", x"6a89",
        x"6a8d", x"6a91", x"6a94", x"6a98", x"6a9c", x"6a9f", x"6aa3", x"6aa7", x"6aab", x"6aae", x"6ab2", x"6ab5", x"6ab9", x"6abd", x"6ac0", x"6ac4",
        x"6ac8", x"6acb", x"6acf", x"6ad2", x"6ad6", x"6ad9", x"6add", x"6ae1", x"6ae4", x"6ae8", x"6aeb", x"6aef", x"6af2", x"6af6", x"6af9", x"6afc",
        x"6b00", x"6b03", x"6b07", x"6b0a", x"6b0e", x"6b11", x"6b14", x"6b18", x"6b1b", x"6b1f", x"6b22", x"6b25", x"6b29", x"6b2c", x"6b2f", x"6b33",
        x"6b36", x"6b39", x"6b3d", x"6b40", x"6b43", x"6b46", x"6b4a", x"6b4d", x"6b50", x"6b53", x"6b57", x"6b5a", x"6b5d", x"6b60", x"6b63", x"6b67",
        x"6b6a", x"6b6d", x"6b70", x"6b73", x"6b76", x"6b7a", x"6b7d", x"6b80", x"6b83", x"6b86", x"6b89", x"6b8c", x"6b8f", x"6b92", x"6b95", x"6b98",
        x"6b9b", x"6b9e", x"6ba1", x"6ba4", x"6ba7", x"6baa", x"6bad", x"6bb0", x"6bb3", x"6bb6", x"6bb9", x"6bbc", x"6bbf", x"6bc2", x"6bc5", x"6bc8",
        x"6bcb", x"6bce", x"6bd1", x"6bd4", x"6bd6", x"6bd9", x"6bdc", x"6bdf", x"6be2", x"6be5", x"6be7", x"6bea", x"6bed", x"6bf0", x"6bf3", x"6bf5",
        x"6bf8", x"6bfb", x"6bfe", x"6c01", x"6c03", x"6c06", x"6c09", x"6c0b", x"6c0e", x"6c11", x"6c14", x"6c16", x"6c19", x"6c1c", x"6c1e", x"6c21",
        x"6c24", x"6c26", x"6c29", x"6c2b", x"6c2e", x"6c31", x"6c33", x"6c36", x"6c39", x"6c3b", x"6c3e", x"6c40", x"6c43", x"6c45", x"6c48", x"6c4a",
        x"6c4d", x"6c4f", x"6c52", x"6c54", x"6c57", x"6c59", x"6c5c", x"6c5e", x"6c61", x"6c63", x"6c66", x"6c68", x"6c6b", x"6c6d", x"6c70", x"6c72",
        x"6c74", x"6c77", x"6c79", x"6c7c", x"6c7e", x"6c80", x"6c83", x"6c85", x"6c87", x"6c8a", x"6c8c", x"6c8e", x"6c91", x"6c93", x"6c95", x"6c98",
        x"6c9a", x"6c9c", x"6c9e", x"6ca1", x"6ca3", x"6ca5", x"6ca7", x"6caa", x"6cac", x"6cae", x"6cb0", x"6cb3", x"6cb5", x"6cb7", x"6cb9", x"6cbb",
        x"6cbe", x"6cc0", x"6cc2", x"6cc4", x"6cc6", x"6cc8", x"6ccb", x"6ccd", x"6ccf", x"6cd1", x"6cd3", x"6cd5", x"6cd7", x"6cd9", x"6cdb", x"6cdd",
        x"6ce0", x"6ce2", x"6ce4", x"6ce6", x"6ce8", x"6cea", x"6cec", x"6cee", x"6cf0", x"6cf2", x"6cf4", x"6cf6", x"6cf8", x"6cfa", x"6cfc", x"6cfe",
        x"6d00", x"6d02", x"6d04", x"6d06", x"6d07", x"6d09", x"6d0b", x"6d0d", x"6d0f", x"6d11", x"6d13", x"6d15", x"6d17", x"6d19", x"6d1a", x"6d1c",
        x"6d1e", x"6d20", x"6d22", x"6d24", x"6d26", x"6d27", x"6d29", x"6d2b", x"6d2d", x"6d2f", x"6d30", x"6d32", x"6d34", x"6d36", x"6d37", x"6d39",
        x"6d3b", x"6d3d", x"6d3e", x"6d40", x"6d42", x"6d44", x"6d45", x"6d47", x"6d49", x"6d4b", x"6d4c", x"6d4e", x"6d50", x"6d51", x"6d53", x"6d55",
        x"6d56", x"6d58", x"6d5a", x"6d5b", x"6d5d", x"6d5e", x"6d60", x"6d62", x"6d63", x"6d65", x"6d66", x"6d68", x"6d6a", x"6d6b", x"6d6d", x"6d6e",
        x"6d70", x"6d72", x"6d73", x"6d75", x"6d76", x"6d78", x"6d79", x"6d7b", x"6d7c", x"6d7e", x"6d7f", x"6d81", x"6d82", x"6d84", x"6d85", x"6d87",
        x"6d88", x"6d8a", x"6d8b", x"6d8d", x"6d8e", x"6d8f", x"6d91", x"6d92", x"6d94", x"6d95", x"6d97", x"6d98", x"6d99", x"6d9b", x"6d9c", x"6d9e",
        x"6d9f", x"6da0", x"6da2", x"6da3", x"6da4", x"6da6", x"6da7", x"6da8", x"6daa", x"6dab", x"6dac", x"6dae", x"6daf", x"6db0", x"6db2", x"6db3",
        x"6db4", x"6db6", x"6db7", x"6db8", x"6db9", x"6dbb", x"6dbc", x"6dbd", x"6dbe", x"6dc0", x"6dc1", x"6dc2", x"6dc3", x"6dc5", x"6dc6", x"6dc7",
        x"6dc8", x"6dc9", x"6dcb", x"6dcc", x"6dcd", x"6dce", x"6dcf", x"6dd1", x"6dd2", x"6dd3", x"6dd4", x"6dd5", x"6dd6", x"6dd8", x"6dd9", x"6dda",
        x"6ddb", x"6ddc", x"6ddd", x"6dde", x"6ddf", x"6de1", x"6de2", x"6de3", x"6de4", x"6de5", x"6de6", x"6de7", x"6de8", x"6de9", x"6dea", x"6deb",
        x"6dec", x"6ded", x"6dee", x"6df0", x"6df1", x"6df2", x"6df3", x"6df4", x"6df5", x"6df6", x"6df7", x"6df8", x"6df9", x"6dfa", x"6dfb", x"6dfc",
        x"6dfd", x"6dfe", x"6dff", x"6e00", x"6e00", x"6e01", x"6e02", x"6e03", x"6e04", x"6e05", x"6e06", x"6e07", x"6e08", x"6e09", x"6e0a", x"6e0b",
        x"6e0c", x"6e0d", x"6e0d", x"6e0e", x"6e0f", x"6e10", x"6e11", x"6e12", x"6e13", x"6e14", x"6e14", x"6e15", x"6e16", x"6e17", x"6e18", x"6e19",
        x"6e1a", x"6e1a", x"6e1b", x"6e1c", x"6e1d", x"6e1e", x"6e1e", x"6e1f", x"6e20", x"6e21", x"6e22", x"6e22", x"6e23", x"6e24", x"6e25", x"6e26",
        x"6e26", x"6e27", x"6e28", x"6e29", x"6e29", x"6e2a", x"6e2b", x"6e2c", x"6e2c", x"6e2d", x"6e2e", x"6e2e", x"6e2f", x"6e30", x"6e31", x"6e31",
        x"6e32", x"6e33", x"6e33", x"6e34", x"6e35", x"6e35", x"6e36", x"6e37", x"6e38", x"6e38", x"6e39", x"6e39", x"6e3a", x"6e3b", x"6e3b", x"6e3c",
        x"6e3d", x"6e3d", x"6e3e", x"6e3f", x"6e3f", x"6e40", x"6e41", x"6e41", x"6e42", x"6e42", x"6e43", x"6e44", x"6e44", x"6e45", x"6e45", x"6e46",
        x"6e46", x"6e47", x"6e48", x"6e48", x"6e49", x"6e49", x"6e4a", x"6e4a", x"6e4b", x"6e4c", x"6e4c", x"6e4d", x"6e4d", x"6e4e", x"6e4e", x"6e4f",
        x"6e4f", x"6e50", x"6e50", x"6e51", x"6e51", x"6e52", x"6e52", x"6e53", x"6e53", x"6e54", x"6e54", x"6e55", x"6e55", x"6e56", x"6e56", x"6e57",
        x"6e57", x"6e58", x"6e58", x"6e59", x"6e59", x"6e59", x"6e5a", x"6e5a", x"6e5b", x"6e5b", x"6e5c", x"6e5c", x"6e5d", x"6e5d", x"6e5d", x"6e5e",
        x"6e5e", x"6e5f", x"6e5f", x"6e5f", x"6e60", x"6e60", x"6e61", x"6e61", x"6e61", x"6e62", x"6e62", x"6e63", x"6e63", x"6e63", x"6e64", x"6e64",
        x"6e64", x"6e65", x"6e65", x"6e66", x"6e66", x"6e66", x"6e67", x"6e67", x"6e67", x"6e68", x"6e68", x"6e68", x"6e69", x"6e69", x"6e69", x"6e6a",
        x"6e6a", x"6e6a", x"6e6b", x"6e6b", x"6e6b", x"6e6b", x"6e6c", x"6e6c", x"6e6c", x"6e6d", x"6e6d", x"6e6d", x"6e6e", x"6e6e", x"6e6e", x"6e6e",
        x"6e6f", x"6e6f", x"6e6f", x"6e6f", x"6e70", x"6e70", x"6e70", x"6e70", x"6e71", x"6e71", x"6e71", x"6e71", x"6e72", x"6e72", x"6e72", x"6e72",
        x"6e73", x"6e73", x"6e73", x"6e73", x"6e74", x"6e74", x"6e74", x"6e74", x"6e74", x"6e75", x"6e75", x"6e75", x"6e75", x"6e75", x"6e76", x"6e76",
        x"6e76", x"6e76", x"6e76", x"6e76", x"6e77", x"6e77", x"6e77", x"6e77", x"6e77", x"6e77", x"6e78", x"6e78", x"6e78", x"6e78", x"6e78", x"6e78",
        x"6e79", x"6e79", x"6e79", x"6e79", x"6e79", x"6e79", x"6e79", x"6e7a", x"6e7a", x"6e7a", x"6e7a", x"6e7a", x"6e7a", x"6e7a", x"6e7a", x"6e7b",
        x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c",
        x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d",
        x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d",
        x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d",
        x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d", x"6e7d",
        x"6e7d", x"6e7d", x"6e7d", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c", x"6e7c",
        x"6e7c", x"6e7c", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7b", x"6e7a", x"6e7a", x"6e7a",
        x"6e7a", x"6e7a", x"6e7a", x"6e7a", x"6e7a", x"6e7a", x"6e7a", x"6e79", x"6e79", x"6e79", x"6e79", x"6e79", x"6e79", x"6e79", x"6e79", x"6e78",
        x"6e78", x"6e78", x"6e78", x"6e78", x"6e78", x"6e78", x"6e78", x"6e77", x"6e77", x"6e77", x"6e77", x"6e77", x"6e77", x"6e77", x"6e76", x"6e76",
        x"6e76", x"6e76", x"6e76", x"6e76", x"6e76", x"6e75", x"6e75", x"6e75", x"6e75", x"6e75", x"6e75", x"6e74", x"6e74", x"6e74", x"6e74", x"6e74",
        x"6e74", x"6e73", x"6e73", x"6e73", x"6e73", x"6e73", x"6e73", x"6e72", x"6e72", x"6e72", x"6e72", x"6e72", x"6e72", x"6e71", x"6e71", x"6e71",
        x"6e71", x"6e71", x"6e70", x"6e70", x"6e70", x"6e70", x"6e70", x"6e6f", x"6e6f", x"6e6f", x"6e6f", x"6e6f", x"6e6e", x"6e6e", x"6e6e", x"6e6e",
        x"6e6e", x"6e6d", x"6e6d", x"6e6d", x"6e6d", x"6e6d", x"6e6c", x"6e6c", x"6e6c", x"6e6c", x"6e6c", x"6e6b", x"6e6b", x"6e6b", x"6e6b", x"6e6a",
        x"6e6a", x"6e6a", x"6e6a", x"6e6a", x"6e69", x"6e69", x"6e69", x"6e69", x"6e68", x"6e68", x"6e68", x"6e68", x"6e68", x"6e67", x"6e67", x"6e67",
        x"6e67", x"6e66", x"6e66", x"6e66", x"6e66", x"6e65", x"6e65", x"6e65", x"6e65", x"6e64", x"6e64", x"6e64", x"6e64", x"6e63", x"6e63", x"6e63",
        x"6e63", x"6e63", x"6e62", x"6e62", x"6e62", x"6e62", x"6e61", x"6e61", x"6e61", x"6e60", x"6e60", x"6e60", x"6e60", x"6e5f", x"6e5f", x"6e5f",
        x"6e5f", x"6e5e", x"6e5e", x"6e5e", x"6e5e", x"6e5d", x"6e5d", x"6e5d", x"6e5d", x"6e5c", x"6e5c", x"6e5c", x"6e5b", x"6e5b", x"6e5b", x"6e5b",
        x"6e5a", x"6e5a", x"6e5a", x"6e5a", x"6e59", x"6e59", x"6e59", x"6e58", x"6e58", x"6e58", x"6e58", x"6e57", x"6e57", x"6e57", x"6e57", x"6e56",
        x"6e56", x"6e56", x"6e55", x"6e55", x"6e55", x"6e55", x"6e54", x"6e54", x"6e54", x"6e53", x"6e53", x"6e53", x"6e53", x"6e52", x"6e52", x"6e52",
        x"6e51", x"6e51", x"6e51", x"6e50", x"6e50", x"6e50", x"6e50", x"6e4f", x"6e4f", x"6e4f", x"6e4e", x"6e4e", x"6e4e", x"6e4e", x"6e4d", x"6e4d",
        x"6e4d", x"6e4c", x"6e4c", x"6e4c", x"6e4b", x"6e4b", x"6e4b", x"6e4b", x"6e4a", x"6e4a", x"6e4a", x"6e49", x"6e49", x"6e49", x"6e48", x"6e48",
        x"6e48", x"6e47", x"6e47", x"6e47", x"6e47", x"6e46", x"6e46", x"6e46", x"6e45", x"6e45", x"6e45", x"6e44", x"6e44", x"6e44", x"6e43", x"6e43",
        x"6e43", x"6e43", x"6e42", x"6e42", x"6e42", x"6e41", x"6e41", x"6e41", x"6e40", x"6e40", x"6e40", x"6e3f", x"6e3f", x"6e3f", x"6e3e", x"6e3e",
        x"6e3e", x"6e3d", x"6e3d", x"6e3d", x"6e3d", x"6e3c", x"6e3c", x"6e3c", x"6e3b", x"6e3b", x"6e3b", x"6e3a", x"6e3a", x"6e3a", x"6e39", x"6e39",
        x"6e39", x"6e38", x"6e38", x"6e38", x"6e37", x"6e37", x"6e37", x"6e36", x"6e36", x"6e36", x"6e35", x"6e35", x"6e35", x"6e34", x"6e34", x"6e34",
        x"6e34", x"6e33", x"6e33", x"6e33", x"6e32", x"6e32", x"6e32", x"6e31", x"6e31", x"6e31", x"6e30", x"6e30", x"6e30", x"6e2f", x"6e2f", x"6e2f",
        x"6e2e", x"6e2e", x"6e2e", x"6e2d", x"6e2d", x"6e2d", x"6e2c", x"6e2c", x"6e2c", x"6e2b", x"6e2b", x"6e2b", x"6e2a", x"6e2a", x"6e2a", x"6e29",
        x"6e29", x"6e29", x"6e28", x"6e28", x"6e28", x"6e27", x"6e27", x"6e27", x"6e26", x"6e26", x"6e26", x"6e25", x"6e25", x"6e25", x"6e24", x"6e24",
        x"6e24", x"6e23", x"6e23", x"6e23", x"6e22", x"6e22", x"6e22", x"6e21", x"6e21", x"6e21", x"6e20", x"6e20", x"6e20", x"6e1f", x"6e1f", x"6e1f",
        x"6e1e", x"6e1e", x"6e1e", x"6e1d", x"6e1d", x"6e1d", x"6e1c", x"6e1c", x"6e1c", x"6e1b", x"6e1b", x"6e1b", x"6e1a", x"6e1a", x"6e1a", x"6e19",
        x"6e19", x"6e19", x"6e18", x"6e18", x"6e18", x"6e17", x"6e17", x"6e17", x"6e16", x"6e16", x"6e16", x"6e15", x"6e15", x"6e15", x"6e14", x"6e14",
        x"6e14", x"6e13", x"6e13", x"6e13", x"6e12", x"6e12", x"6e12", x"6e11", x"6e11", x"6e11", x"6e10", x"6e10", x"6e10", x"6e10", x"6e0f", x"6e0f",
        x"6e0f", x"6e0e", x"6e0e", x"6e0e", x"6e0d", x"6e0d", x"6e0d", x"6e0c", x"6e0c", x"6e0c", x"6e0b", x"6e0b", x"6e0b", x"6e0a", x"6e0a", x"6e0a",
        x"6e09", x"6e09", x"6e09", x"6e08", x"6e08", x"6e08", x"6e07", x"6e07", x"6e07", x"6e06", x"6e06", x"6e06", x"6e05", x"6e05", x"6e05", x"6e04",
        x"6e04", x"6e04", x"6e03", x"6e03", x"6e03", x"6e02", x"6e02", x"6e02", x"6e01", x"6e01", x"6e01", x"6e00", x"6e00", x"6e00", x"6dff", x"6dff",
        x"6dff", x"6dff", x"6dfe", x"6dfe", x"6dfe", x"6dfd", x"6dfd", x"6dfd", x"6dfc", x"6dfc", x"6dfc", x"6dfb", x"6dfb", x"6dfb", x"6dfa", x"6dfa",
        x"6dfa", x"6df9", x"6df9", x"6df9", x"6df8", x"6df8", x"6df8", x"6df7", x"6df7", x"6df7", x"6df6", x"6df6", x"6df6", x"6df6", x"6df5", x"6df5",
        x"6df5", x"6df4", x"6df4", x"6df4", x"6df3", x"6df3", x"6df3", x"6df2", x"6df2", x"6df2", x"6df1", x"6df1", x"6df1", x"6df0", x"6df0", x"6df0",
        x"6df0", x"6def", x"6def", x"6def", x"6dee", x"6dee", x"6dee", x"6ded", x"6ded", x"6ded", x"6dec", x"6dec", x"6dec", x"6dec", x"6deb", x"6deb",
        x"6deb", x"6dea", x"6dea", x"6dea", x"6de9", x"6de9", x"6de9", x"6de8", x"6de8", x"6de8", x"6de8", x"6de7", x"6de7", x"6de7", x"6de6", x"6de6",
        x"6de6", x"6de5", x"6de5", x"6de5", x"6de4", x"6de4", x"6de4", x"6de4", x"6de3", x"6de3", x"6de3", x"6de2", x"6de2", x"6de2", x"6de1", x"6de1",
        x"6de1", x"6de1", x"6de0", x"6de0", x"6de0", x"6ddf", x"6ddf", x"6ddf", x"6dde", x"6dde", x"6dde", x"6dde", x"6ddd", x"6ddd", x"6ddd", x"6ddc",
        x"6ddc", x"6ddc", x"6ddc", x"6ddb", x"6ddb", x"6ddb", x"6dda", x"6dda", x"6dda", x"6dda", x"6dd9", x"6dd9", x"6dd9", x"6dd8", x"6dd8", x"6dd8",
        x"6dd7", x"6dd7", x"6dd7", x"6dd7", x"6dd6", x"6dd6", x"6dd6", x"6dd5", x"6dd5", x"6dd5", x"6dd5", x"6dd4", x"6dd4", x"6dd4", x"6dd3", x"6dd3",
        x"6dd3", x"6dd3", x"6dd2", x"6dd2", x"6dd2", x"6dd1", x"6dd1", x"6dd1", x"6dd1", x"6dd0", x"6dd0", x"6dd0", x"6dd0", x"6dcf", x"6dcf", x"6dcf",
        x"6dce", x"6dce", x"6dce", x"6dce", x"6dcd", x"6dcd", x"6dcd", x"6dcc", x"6dcc", x"6dcc", x"6dcc", x"6dcb", x"6dcb", x"6dcb", x"6dcb", x"6dca",
        x"6dca", x"6dca", x"6dca", x"6dc9", x"6dc9", x"6dc9", x"6dc8", x"6dc8", x"6dc8", x"6dc8", x"6dc7", x"6dc7", x"6dc7", x"6dc7", x"6dc6", x"6dc6",
        x"6dc6", x"6dc5", x"6dc5", x"6dc5", x"6dc5", x"6dc4", x"6dc4", x"6dc4", x"6dc4", x"6dc3", x"6dc3", x"6dc3", x"6dc3", x"6dc2", x"6dc2", x"6dc2",
        x"6dc2", x"6dc1", x"6dc1", x"6dc1", x"6dc1", x"6dc0", x"6dc0", x"6dc0", x"6dc0", x"6dbf", x"6dbf", x"6dbf", x"6dbe", x"6dbe", x"6dbe", x"6dbe",
        x"6dbd", x"6dbd", x"6dbd", x"6dbd", x"6dbc", x"6dbc", x"6dbc", x"6dbc", x"6dbb", x"6dbb", x"6dbb", x"6dbb", x"6dba", x"6dba", x"6dba", x"6dba",
        x"6db9", x"6db9", x"6db9", x"6db9", x"6db9", x"6db8", x"6db8", x"6db8", x"6db8", x"6db7", x"6db7", x"6db7", x"6db7", x"6db6", x"6db6", x"6db6",
        x"6db6", x"6db5", x"6db5", x"6db5", x"6db5", x"6db4", x"6db4", x"6db4", x"6db4", x"6db3", x"6db3", x"6db3", x"6db3", x"6db3", x"6db2", x"6db2",
        x"6db2", x"6db2", x"6db1", x"6db1", x"6db1", x"6db1", x"6db0", x"6db0", x"6db0", x"6db0", x"6db0", x"6daf", x"6daf", x"6daf", x"6daf", x"6dae",
        x"6dae", x"6dae", x"6dae", x"6dad", x"6dad", x"6dad", x"6dad", x"6dad", x"6dac", x"6dac", x"6dac", x"6dac", x"6dab", x"6dab", x"6dab", x"6dab",
        x"6dab", x"6daa", x"6daa", x"6daa", x"6daa", x"6daa", x"6da9", x"6da9", x"6da9", x"6da9", x"6da8", x"6da8", x"6da8", x"6da8", x"6da8", x"6da7",
        x"6da7", x"6da7", x"6da7", x"6da6", x"6da6", x"6da6", x"6da6", x"6da6", x"6da5", x"6da5", x"6da5", x"6da5", x"6da5", x"6da4", x"6da4", x"6da4",
        x"6da4", x"6da4", x"6da3", x"6da3", x"6da3", x"6da3", x"6da3", x"6da2", x"6da2", x"6da2", x"6da2", x"6da2", x"6da1", x"6da1", x"6da1", x"6da1",
        x"6da1", x"6da0", x"6da0", x"6da0", x"6da0", x"6da0", x"6d9f", x"6d9f", x"6d9f", x"6d9f", x"6d9f", x"6d9e", x"6d9e", x"6d9e", x"6d9e", x"6d9e",
        x"6d9d", x"6d9d", x"6d9d", x"6d9d", x"6d9d", x"6d9c", x"6d9c", x"6d9c", x"6d9c", x"6d9c", x"6d9b", x"6d9b", x"6d9b", x"6d9b", x"6d9b", x"6d9b",
        x"6d9a", x"6d9a", x"6d9a", x"6d9a", x"6d9a", x"6d99", x"6d99", x"6d99", x"6d99", x"6d99", x"6d99", x"6d98", x"6d98", x"6d98", x"6d98", x"6d98",
        x"6d97", x"6d97", x"6d97", x"6d97", x"6d97", x"6d97", x"6d96", x"6d96", x"6d96", x"6d96", x"6d96", x"6d95", x"6d95", x"6d95", x"6d95", x"6d95",
        x"6d95", x"6d94", x"6d94", x"6d94", x"6d94", x"6d94", x"6d94", x"6d93", x"6d93", x"6d93", x"6d93", x"6d93", x"6d93", x"6d92", x"6d92", x"6d92",
        x"6d92", x"6d92", x"6d92", x"6d91", x"6d91", x"6d91", x"6d91", x"6d91", x"6d91", x"6d90", x"6d90", x"6d90", x"6d90", x"6d90", x"6d90", x"6d8f",
        x"6d8f", x"6d8f", x"6d8f", x"6d8f", x"6d8f", x"6d8e", x"6d8e", x"6d8e", x"6d8e", x"6d8e", x"6d8e", x"6d8d", x"6d8d", x"6d8d", x"6d8d", x"6d8d",
        x"6d8d", x"6d8d", x"6d8c", x"6d8c", x"6d8c", x"6d8c", x"6d8c", x"6d8c", x"6d8b", x"6d8b", x"6d8b", x"6d8b", x"6d8b", x"6d8b", x"6d8b", x"6d8a",
        x"6d8a", x"6d8a", x"6d8a", x"6d8a", x"6d8a", x"6d8a", x"6d89", x"6d89", x"6d89", x"6d89", x"6d89", x"6d89", x"6d89", x"6d88", x"6d88", x"6d88",
        x"6d88", x"6d88", x"6d88", x"6d88", x"6d87", x"6d87", x"6d87", x"6d87", x"6d87", x"6d87", x"6d87", x"6d86", x"6d86", x"6d86", x"6d86", x"6d86",
        x"6d86", x"6d86", x"6d85", x"6d85", x"6d85", x"6d85", x"6d85", x"6d85", x"6d85", x"6d84", x"6d84", x"6d84", x"6d84", x"6d84", x"6d84", x"6d84",
        x"6d84", x"6d83", x"6d83", x"6d83", x"6d83", x"6d83", x"6d83", x"6d83", x"6d83", x"6d82", x"6d82", x"6d82", x"6d82", x"6d82", x"6d82", x"6d82",
        x"6d81", x"6d81", x"6d81", x"6d81", x"6d81", x"6d81", x"6d81", x"6d81", x"6d80", x"6d80", x"6d80", x"6d80", x"6d80", x"6d80", x"6d80", x"6d80",
        x"6d80", x"6d7f", x"6d7f", x"6d7f", x"6d7f", x"6d7f", x"6d7f", x"6d7f", x"6d7f", x"6d7e", x"6d7e", x"6d7e", x"6d7e", x"6d7e", x"6d7e", x"6d7e",
        x"6d7e", x"6d7e", x"6d7d", x"6d7d", x"6d7d", x"6d7d", x"6d7d", x"6d7d", x"6d7d", x"6d7d", x"6d7c", x"6d7c", x"6d7c", x"6d7c", x"6d7c", x"6d7c",
        x"6d7c", x"6d7c", x"6d7c", x"6d7b", x"6d7b", x"6d7b", x"6d7b", x"6d7b", x"6d7b", x"6d7b", x"6d7b", x"6d7b", x"6d7b", x"6d7a", x"6d7a", x"6d7a",
        x"6d7a", x"6d7a", x"6d7a", x"6d7a", x"6d7a", x"6d7a", x"6d79", x"6d79", x"6d79", x"6d79", x"6d79", x"6d79", x"6d79", x"6d79", x"6d79", x"6d79",
        x"6d78", x"6d78", x"6d78", x"6d78", x"6d78", x"6d78", x"6d78", x"6d78", x"6d78", x"6d78", x"6d77", x"6d77", x"6d77", x"6d77", x"6d77", x"6d77",
        x"6d77", x"6d77", x"6d77", x"6d77", x"6d77", x"6d76", x"6d76", x"6d76", x"6d76", x"6d76", x"6d76", x"6d76", x"6d76", x"6d76", x"6d76", x"6d75",
        x"6d75", x"6d75", x"6d75", x"6d75", x"6d75", x"6d75", x"6d75", x"6d75", x"6d75", x"6d75", x"6d75", x"6d74", x"6d74", x"6d74", x"6d74", x"6d74",
        x"6d74", x"6d74", x"6d74", x"6d74", x"6d74", x"6d74", x"6d73", x"6d73", x"6d73", x"6d73", x"6d73", x"6d73", x"6d73", x"6d73", x"6d73", x"6d73",
        x"6d73", x"6d73", x"6d72", x"6d72", x"6d72", x"6d72", x"6d72", x"6d72", x"6d72", x"6d72", x"6d72", x"6d72", x"6d72", x"6d72", x"6d71", x"6d71",
        x"6d71", x"6d71", x"6d71", x"6d71", x"6d71", x"6d71", x"6d71", x"6d71", x"6d71", x"6d71", x"6d71", x"6d70", x"6d70", x"6d70", x"6d70", x"6d70",
        x"6d70", x"6d70", x"6d70", x"6d70", x"6d70", x"6d70", x"6d70", x"6d70", x"6d70", x"6d6f", x"6d6f", x"6d6f", x"6d6f", x"6d6f", x"6d6f", x"6d6f",
        x"6d6f", x"6d6f", x"6d6f", x"6d6f", x"6d6f", x"6d6f", x"6d6f", x"6d6e", x"6d6e", x"6d6e", x"6d6e", x"6d6e", x"6d6e", x"6d6e", x"6d6e", x"6d6e",
        x"6d6e", x"6d6e", x"6d6e", x"6d6e", x"6d6e", x"6d6e", x"6d6d", x"6d6d", x"6d6d", x"6d6d", x"6d6d", x"6d6d", x"6d6d", x"6d6d", x"6d6d", x"6d6d",
        x"6d6d", x"6d6d", x"6d6d", x"6d6d", x"6d6d", x"6d6c", x"6d6c", x"6d6c", x"6d6c", x"6d6c", x"6d6c", x"6d6c", x"6d6c", x"6d6c", x"6d6c", x"6d6c",
        x"6d6c", x"6d6c", x"6d6c", x"6d6c", x"6d6c", x"6d6b", x"6d6b", x"6d6b", x"6d6b", x"6d6b", x"6d6b", x"6d6b", x"6d6b", x"6d6b", x"6d6b", x"6d6b",
        x"6d6b", x"6d6b", x"6d6b", x"6d6b", x"6d6b", x"6d6b", x"6d6b", x"6d6a", x"6d6a", x"6d6a", x"6d6a", x"6d6a", x"6d6a", x"6d6a", x"6d6a", x"6d6a",
        x"6d6a", x"6d6a", x"6d6a", x"6d6a", x"6d6a", x"6d6a", x"6d6a", x"6d6a", x"6d6a", x"6d69", x"6d69", x"6d69", x"6d69", x"6d69", x"6d69", x"6d69",
        x"6d69", x"6d69", x"6d69", x"6d69", x"6d69", x"6d69", x"6d69", x"6d69", x"6d69", x"6d69", x"6d69", x"6d69", x"6d68", x"6d68", x"6d68", x"6d68",
        x"6d68", x"6d68", x"6d68", x"6d68", x"6d68", x"6d68", x"6d68", x"6d68", x"6d68", x"6d68", x"6d68", x"6d68", x"6d68", x"6d68", x"6d68", x"6d68",
        x"6d68", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67",
        x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d67", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66",
        x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d66", x"6d65", x"6d65",
        x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65",
        x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d65", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64",
        x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64", x"6d64",
        x"6d64", x"6d64", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63",
        x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d63", x"6d62",
        x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62",
        x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d62", x"6d61", x"6d61",
        x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61",
        x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d61", x"6d60", x"6d60",
        x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60",
        x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60", x"6d60"
           );

   signal state : std_logic_vector(1 downto 0) := "00";
   signal count : unsigned(12 downto 0) := (others => '0');

begin

process(clk)
   begin
      if rising_edge(clk) then
         baseband <= lookup(to_integer(count));
         case state is
            when "00" => 
               if tx = '1' then
                  state <= "01";
               end if;
            when "01" =>
               count <= count + 1;
               if count = 8190 then
                  state <= "10";
               end if;
            when "10" =>
               if tx = '0' then
                  state <= "11";
               end if;
            when "11" =>
               count <= count - 1;
               if count = 1 then
                  state <= "00";
               end if;
            when others =>
               state <= "00";
         end case;
      end if;
   end process;
end Behavioral;
